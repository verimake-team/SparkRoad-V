// Verilog netlist created by TD v4.5.12562
// Mon Sep 30 17:08:52 2019

`timescale 1ns / 1ps
module M0demo  // ../RTL/M0demo.v(4)
  (
  NRST,
  SWCLKTCK,
  TDI,
  XTAL1,
  nTRST,
  uart0_rxd,
  P0,
  TDO,
  XTAL2,
  uart0_txd,
  uart0_txen,
  SWDIOTMS,
  b_pad_gpio_porta
  );

  input NRST;  // ../RTL/M0demo.v(7)
  input SWCLKTCK;  // ../RTL/M0demo.v(15)
  input TDI;  // ../RTL/M0demo.v(12)
  input XTAL1;  // ../RTL/M0demo.v(5)
  input nTRST;  // ../RTL/M0demo.v(11)
  input uart0_rxd;  // ../RTL/M0demo.v(19)
  output [15:0] P0;  // ../RTL/M0demo.v(8)
  output TDO;  // ../RTL/M0demo.v(13)
  output XTAL2;  // ../RTL/M0demo.v(6)
  output uart0_txd;  // ../RTL/M0demo.v(20)
  output uart0_txen;  // ../RTL/M0demo.v(21)
  inout SWDIOTMS;  // ../RTL/M0demo.v(14)
  inout [7:0] b_pad_gpio_porta;  // ../RTL/M0demo.v(17)

  parameter BE = 0;
  parameter BKPT = 4;
  parameter DBG = 1;
  parameter NUMIRQ = 32;
  parameter SMUL = 0;
  parameter SYST = 1;
  parameter WIC = 1;
  parameter WICLINES = 34;
  parameter WPT = 2;
  wire [7:0] b_pad_gpio_porta_pad;  // ../RTL/M0demo.v(17)
  wire [13:0] n0;
  wire [13:0] n1;
  wire [31:0] \u_cmsdk_mcu/HADDR ;  // ../RTL/cmsdk_mcu.v(103)
  wire [2:0] \u_cmsdk_mcu/HSIZE ;  // ../RTL/cmsdk_mcu.v(105)
  wire [1:0] \u_cmsdk_mcu/HTRANS ;  // ../RTL/cmsdk_mcu.v(104)
  wire [31:0] \u_cmsdk_mcu/HWDATA ;  // ../RTL/cmsdk_mcu.v(107)
  wire [31:0] \u_cmsdk_mcu/flash_hrdata ;  // ../RTL/cmsdk_mcu.v(113)
  wire [15:0] \u_cmsdk_mcu/p0_altfunc ;  // ../RTL/cmsdk_mcu.v(140)
  wire [15:0] \u_cmsdk_mcu/p0_out ;  // ../RTL/cmsdk_mcu.v(138)
  wire [15:0] \u_cmsdk_mcu/p0_outen ;  // ../RTL/cmsdk_mcu.v(139)
  wire [15:0] \u_cmsdk_mcu/p1_altfunc ;  // ../RTL/cmsdk_mcu.v(145)
  wire [15:0] \u_cmsdk_mcu/p1_out ;  // ../RTL/cmsdk_mcu.v(143)
  wire [15:0] \u_cmsdk_mcu/p1_outen ;  // ../RTL/cmsdk_mcu.v(144)
  wire [31:0] \u_cmsdk_mcu/sram_hrdata ;  // ../RTL/cmsdk_mcu.v(119)
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/buf_hwaddr ;  // ../RTL/AHB2MEM.v(30)
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/hwdata_mask ;  // ../RTL/AHB2MEM.v(28)
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/n13 ;
  wire [31:0] \u_cmsdk_mcu/u_ahb_ram/n5 ;
  wire [31:0] \u_cmsdk_mcu/u_ahb_rom/n13 ;
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg ;  // ../RTL/cmsdk_mcu_clkctrl.v(62)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt ;  // ../RTL/cmsdk_mcu_system.v(307)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr ;  // ../RTL/cmsdk_mcu_system.v(304)
  wire [11:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR ;  // ../RTL/cmsdk_ahb_gpio.v(76)
  wire [1:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE ;  // ../RTL/cmsdk_ahb_gpio.v(78)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 ;
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int ;  // ../RTL/cmsdk_iop_gpio.v(517)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded ;  // ../RTL/cmsdk_iop_gpio.v(397)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded ;  // ../RTL/cmsdk_iop_gpio.v(474)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded ;  // ../RTL/cmsdk_iop_gpio.v(435)
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b0/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b1/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b10/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b11/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b12/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b13/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b14/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b15/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b2/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b3/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b4/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b5/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b6/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b7/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b8/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b9/B1_0 ;
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int ;  // ../RTL/cmsdk_iop_gpio.v(517)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int ;  // ../RTL/cmsdk_iop_gpio.v(129)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 ;  // ../RTL/cmsdk_iop_gpio.v(238)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 ;  // ../RTL/cmsdk_iop_gpio.v(239)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded ;  // ../RTL/cmsdk_iop_gpio.v(397)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded ;  // ../RTL/cmsdk_iop_gpio.v(474)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded ;  // ../RTL/cmsdk_iop_gpio.v(435)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain ;  // ../RTL/cmsdk_iop_gpio.v(549)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n35 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 ;
  wire [9:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel ;  // ../RTL/cmsdk_ahb_slave_mux.v(95)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity ;  // ../RTL/gpio.v(60)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten ;  // ../RTL/gpio.v(61)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask ;  // ../RTL/gpio.v(62)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level ;  // ../RTL/gpio.v(67)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus ;  // ../RTL/gpio.v(73)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr ;  // ../RTL/gpio.v(75)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr ;  // ../RTL/gpio.v(76)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync ;  // ../RTL/gpio_apbif.v(98)
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b0/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b1/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b2/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b3/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b4/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b5/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b6/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b7/B1_0 ;
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 ;  // ../RTL/gpio_ctrl.v(70)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int ;  // ../RTL/gpio_ctrl.v(72)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm ;  // ../RTL/gpio_ctrl.v(74)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in ;  // ../RTL/gpio_ctrl.v(79)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 ;  // ../RTL/gpio_ctrl.v(80)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in ;  // ../RTL/gpio_ctrl.v(83)
  wire [1:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set ;  // ../RTL/cmsdk_apb_uart.v(147)
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b4/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b5/B1_0 ;
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b6/B1_0 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 ;
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n26 ;
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 ;
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 ;
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 ;
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg ;  // ../RTL/cmsdk_apb_uart.v(110)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f ;  // ../RTL/cmsdk_apb_uart.v(124)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i ;  // ../RTL/cmsdk_apb_uart.v(122)
  wire [19:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div ;  // ../RTL/cmsdk_apb_uart.v(118)
  wire [6:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl ;  // ../RTL/cmsdk_apb_uart.v(115)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf ;  // ../RTL/cmsdk_apb_uart.v(117)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf ;  // ../RTL/cmsdk_apb_uart.v(116)
  wire [6:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf ;  // ../RTL/cmsdk_apb_uart.v(182)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state ;  // ../RTL/cmsdk_apb_uart.v(175)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(178)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf ;  // ../RTL/cmsdk_apb_uart.v(170)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf ;  // ../RTL/cmsdk_apb_uart.v(157)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state ;  // ../RTL/cmsdk_apb_uart.v(151)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(155)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(185)
  wire [15:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(170)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg ;  // ../RTL/cmsdk_ahb_to_apb.v(90)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg ;  // ../RTL/cmsdk_ahb_to_apb.v(80)
  wire  \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux3_b0/B1_0 ;
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 ;
  wire [11:2] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr ;  // ../RTL/cmsdk_mcu_sysctrl.v(123)
  wire [3:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe ;  // ../RTL/cmsdk_mcu_sysctrl.v(120)
  wire [2:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo ;  // ../RTL/cmsdk_mcu_sysctrl.v(109)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 ;  // ../RTL/cortexm0ds_logic.v(1528)
  wire [23:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 ;  // ../RTL/cortexm0ds_logic.v(1545)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 ;  // ../RTL/cortexm0ds_logic.v(1531)
  wire [30:2] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 ;  // ../RTL/cortexm0ds_logic.v(1523)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 ;  // ../RTL/cortexm0ds_logic.v(1719)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 ;  // ../RTL/cortexm0ds_logic.v(1720)
  wire [33:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 ;  // ../RTL/cortexm0ds_logic.v(1721)
  wire [30:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 ;  // ../RTL/cortexm0ds_logic.v(1527)
  wire [31:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 ;  // ../RTL/cortexm0ds_logic.v(1530)
  wire [7:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 ;  // ../RTL/cortexm0ds_logic.v(1534)
  wire [33:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 ;  // ../RTL/cortexm0ds_logic.v(1718)
  wire [8:1] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 ;  // ../RTL/cortexm0ds_logic.v(1533)
  wire [30:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 ;  // ../RTL/cortexm0ds_logic.v(1537)
  wire [9:0] \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg ;  // ../RTL/cmsdk_ahb_cs_rom_table.v(118)
  wire NRST_pad;  // ../RTL/M0demo.v(7)
  wire SWCLKTCK_pad;  // ../RTL/M0demo.v(15)
  wire XTAL1_pad;  // ../RTL/M0demo.v(5)
  wire XTAL1_wire;  // ../RTL/M0demo.v(25)
  wire XTAL2_pad;  // ../RTL/M0demo.v(6)
  wire _al_u1000_o;
  wire _al_u1001_o;
  wire _al_u1002_o;
  wire _al_u1003_o;
  wire _al_u1004_o;
  wire _al_u1006_o;
  wire _al_u1008_o;
  wire _al_u1010_o;
  wire _al_u1011_o;
  wire _al_u1012_o;
  wire _al_u1013_o;
  wire _al_u1015_o;
  wire _al_u1016_o;
  wire _al_u1017_o;
  wire _al_u1018_o;
  wire _al_u1020_o;
  wire _al_u1023_o;
  wire _al_u1024_o;
  wire _al_u1025_o;
  wire _al_u1026_o;
  wire _al_u1027_o;
  wire _al_u1028_o;
  wire _al_u1030_o;
  wire _al_u1032_o;
  wire _al_u1033_o;
  wire _al_u1034_o;
  wire _al_u1035_o;
  wire _al_u1039_o;
  wire _al_u1040_o;
  wire _al_u1048_o;
  wire _al_u1055_o;
  wire _al_u1058_o;
  wire _al_u1061_o;
  wire _al_u1064_o;
  wire _al_u1065_o;
  wire _al_u1066_o;
  wire _al_u1070_o;
  wire _al_u1071_o;
  wire _al_u1073_o;
  wire _al_u1076_o;
  wire _al_u1077_o;
  wire _al_u1078_o;
  wire _al_u1079_o;
  wire _al_u1082_o;
  wire _al_u1083_o;
  wire _al_u1085_o;
  wire _al_u1088_o;
  wire _al_u1089_o;
  wire _al_u1090_o;
  wire _al_u1091_o;
  wire _al_u1094_o;
  wire _al_u1095_o;
  wire _al_u1096_o;
  wire _al_u1097_o;
  wire _al_u1100_o;
  wire _al_u1101_o;
  wire _al_u1102_o;
  wire _al_u1103_o;
  wire _al_u1106_o;
  wire _al_u1107_o;
  wire _al_u1109_o;
  wire _al_u1112_o;
  wire _al_u1113_o;
  wire _al_u1114_o;
  wire _al_u1115_o;
  wire _al_u1118_o;
  wire _al_u1119_o;
  wire _al_u1121_o;
  wire _al_u1124_o;
  wire _al_u1125_o;
  wire _al_u1126_o;
  wire _al_u1131_o;
  wire _al_u1132_o;
  wire _al_u1133_o;
  wire _al_u1137_o;
  wire _al_u1138_o;
  wire _al_u1139_o;
  wire _al_u1142_o;
  wire _al_u1143_o;
  wire _al_u1144_o;
  wire _al_u1145_o;
  wire _al_u1148_o;
  wire _al_u1149_o;
  wire _al_u1150_o;
  wire _al_u1151_o;
  wire _al_u1154_o;
  wire _al_u1155_o;
  wire _al_u1156_o;
  wire _al_u1157_o;
  wire _al_u1160_o;
  wire _al_u1161_o;
  wire _al_u1162_o;
  wire _al_u1163_o;
  wire _al_u1166_o;
  wire _al_u1167_o;
  wire _al_u1168_o;
  wire _al_u1169_o;
  wire _al_u1173_o;
  wire _al_u1174_o;
  wire _al_u1175_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u1181_o;
  wire _al_u1184_o;
  wire _al_u1185_o;
  wire _al_u1186_o;
  wire _al_u1187_o;
  wire _al_u1190_o;
  wire _al_u1193_o;
  wire _al_u1196_o;
  wire _al_u1197_o;
  wire _al_u1198_o;
  wire _al_u1202_o;
  wire _al_u1203_o;
  wire _al_u1204_o;
  wire _al_u1208_o;
  wire _al_u1209_o;
  wire _al_u1210_o;
  wire _al_u1211_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1217_o;
  wire _al_u1220_o;
  wire _al_u1221_o;
  wire _al_u1223_o;
  wire _al_u1226_o;
  wire _al_u1227_o;
  wire _al_u1228_o;
  wire _al_u1229_o;
  wire _al_u1232_o;
  wire _al_u1233_o;
  wire _al_u1234_o;
  wire _al_u1235_o;
  wire _al_u1238_o;
  wire _al_u1239_o;
  wire _al_u1240_o;
  wire _al_u1241_o;
  wire _al_u1244_o;
  wire _al_u1245_o;
  wire _al_u1246_o;
  wire _al_u1247_o;
  wire _al_u1250_o;
  wire _al_u1251_o;
  wire _al_u1253_o;
  wire _al_u1255_o;
  wire _al_u1257_o;
  wire _al_u1264_o;
  wire _al_u1266_o;
  wire _al_u1268_o;
  wire _al_u1269_o;
  wire _al_u1270_o;
  wire _al_u1271_o;
  wire _al_u1273_o;
  wire _al_u1276_o;
  wire _al_u1281_o;
  wire _al_u1282_o;
  wire _al_u1285_o;
  wire _al_u1286_o;
  wire _al_u1288_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1296_o;
  wire _al_u1297_o;
  wire _al_u1299_o;
  wire _al_u1301_o;
  wire _al_u1304_o;
  wire _al_u1305_o;
  wire _al_u1307_o;
  wire _al_u1308_o;
  wire _al_u1309_o;
  wire _al_u1310_o;
  wire _al_u1311_o;
  wire _al_u1316_o;
  wire _al_u1319_o;
  wire _al_u1323_o;
  wire _al_u1327_o;
  wire _al_u1328_o;
  wire _al_u1329_o;
  wire _al_u1331_o;
  wire _al_u1332_o;
  wire _al_u1333_o;
  wire _al_u1334_o;
  wire _al_u1336_o;
  wire _al_u1337_o;
  wire _al_u1339_o;
  wire _al_u1341_o;
  wire _al_u1342_o;
  wire _al_u1343_o;
  wire _al_u1344_o;
  wire _al_u1345_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1354_o;
  wire _al_u1357_o;
  wire _al_u1359_o;
  wire _al_u1360_o;
  wire _al_u1363_o;
  wire _al_u1364_o;
  wire _al_u1366_o;
  wire _al_u1367_o;
  wire _al_u1370_o;
  wire _al_u1372_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1379_o;
  wire _al_u1380_o;
  wire _al_u1381_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1385_o;
  wire _al_u1387_o;
  wire _al_u1390_o;
  wire _al_u1391_o;
  wire _al_u1393_o;
  wire _al_u1394_o;
  wire _al_u1395_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1399_o;
  wire _al_u1400_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1403_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1409_o;
  wire _al_u1410_o;
  wire _al_u1411_o;
  wire _al_u1412_o;
  wire _al_u1413_o;
  wire _al_u1415_o;
  wire _al_u1416_o;
  wire _al_u1417_o;
  wire _al_u1418_o;
  wire _al_u1419_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1423_o;
  wire _al_u1424_o;
  wire _al_u1425_o;
  wire _al_u1426_o;
  wire _al_u1427_o;
  wire _al_u1428_o;
  wire _al_u1429_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1433_o;
  wire _al_u1435_o;
  wire _al_u1436_o;
  wire _al_u1437_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1441_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1445_o;
  wire _al_u1447_o;
  wire _al_u1448_o;
  wire _al_u1449_o;
  wire _al_u1450_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1453_o;
  wire _al_u1455_o;
  wire _al_u1456_o;
  wire _al_u1457_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1460_o;
  wire _al_u1461_o;
  wire _al_u1463_o;
  wire _al_u1464_o;
  wire _al_u1465_o;
  wire _al_u1466_o;
  wire _al_u1467_o;
  wire _al_u1468_o;
  wire _al_u1469_o;
  wire _al_u1471_o;
  wire _al_u1472_o;
  wire _al_u1473_o;
  wire _al_u1474_o;
  wire _al_u1475_o;
  wire _al_u1476_o;
  wire _al_u1477_o;
  wire _al_u1479_o;
  wire _al_u1480_o;
  wire _al_u1481_o;
  wire _al_u1483_o;
  wire _al_u1484_o;
  wire _al_u1485_o;
  wire _al_u1487_o;
  wire _al_u1488_o;
  wire _al_u1489_o;
  wire _al_u1490_o;
  wire _al_u1491_o;
  wire _al_u1492_o;
  wire _al_u1493_o;
  wire _al_u1495_o;
  wire _al_u1496_o;
  wire _al_u1497_o;
  wire _al_u1498_o;
  wire _al_u1499_o;
  wire _al_u1500_o;
  wire _al_u1503_o;
  wire _al_u1504_o;
  wire _al_u1505_o;
  wire _al_u1506_o;
  wire _al_u1507_o;
  wire _al_u1508_o;
  wire _al_u1511_o;
  wire _al_u1512_o;
  wire _al_u1513_o;
  wire _al_u1514_o;
  wire _al_u1515_o;
  wire _al_u1516_o;
  wire _al_u1519_o;
  wire _al_u1520_o;
  wire _al_u1521_o;
  wire _al_u1522_o;
  wire _al_u1523_o;
  wire _al_u1524_o;
  wire _al_u1525_o;
  wire _al_u1527_o;
  wire _al_u1528_o;
  wire _al_u1529_o;
  wire _al_u1531_o;
  wire _al_u1532_o;
  wire _al_u1533_o;
  wire _al_u1535_o;
  wire _al_u1536_o;
  wire _al_u1537_o;
  wire _al_u1538_o;
  wire _al_u1539_o;
  wire _al_u1540_o;
  wire _al_u1541_o;
  wire _al_u1543_o;
  wire _al_u1544_o;
  wire _al_u1545_o;
  wire _al_u1546_o;
  wire _al_u1547_o;
  wire _al_u1548_o;
  wire _al_u1551_o;
  wire _al_u1552_o;
  wire _al_u1553_o;
  wire _al_u1554_o;
  wire _al_u1555_o;
  wire _al_u1556_o;
  wire _al_u1559_o;
  wire _al_u1560_o;
  wire _al_u1561_o;
  wire _al_u1562_o;
  wire _al_u1563_o;
  wire _al_u1564_o;
  wire _al_u1567_o;
  wire _al_u1568_o;
  wire _al_u1569_o;
  wire _al_u1570_o;
  wire _al_u1571_o;
  wire _al_u1572_o;
  wire _al_u1573_o;
  wire _al_u1575_o;
  wire _al_u1576_o;
  wire _al_u1577_o;
  wire _al_u1578_o;
  wire _al_u1579_o;
  wire _al_u1580_o;
  wire _al_u1581_o;
  wire _al_u1582_o;
  wire _al_u1583_o;
  wire _al_u1584_o;
  wire _al_u1586_o;
  wire _al_u1587_o;
  wire _al_u1588_o;
  wire _al_u1589_o;
  wire _al_u1590_o;
  wire _al_u1591_o;
  wire _al_u1592_o;
  wire _al_u1594_o;
  wire _al_u1595_o;
  wire _al_u1596_o;
  wire _al_u1597_o;
  wire _al_u1598_o;
  wire _al_u1599_o;
  wire _al_u1600_o;
  wire _al_u1602_o;
  wire _al_u1603_o;
  wire _al_u1604_o;
  wire _al_u1605_o;
  wire _al_u1606_o;
  wire _al_u1607_o;
  wire _al_u1608_o;
  wire _al_u1610_o;
  wire _al_u1611_o;
  wire _al_u1612_o;
  wire _al_u1613_o;
  wire _al_u1614_o;
  wire _al_u1615_o;
  wire _al_u1616_o;
  wire _al_u1618_o;
  wire _al_u1619_o;
  wire _al_u1620_o;
  wire _al_u1621_o;
  wire _al_u1622_o;
  wire _al_u1623_o;
  wire _al_u1624_o;
  wire _al_u1626_o;
  wire _al_u1627_o;
  wire _al_u1628_o;
  wire _al_u1629_o;
  wire _al_u1630_o;
  wire _al_u1631_o;
  wire _al_u1632_o;
  wire _al_u1634_o;
  wire _al_u1635_o;
  wire _al_u1636_o;
  wire _al_u1638_o;
  wire _al_u1642_o;
  wire _al_u1643_o;
  wire _al_u1644_o;
  wire _al_u1646_o;
  wire _al_u1648_o;
  wire _al_u1652_o;
  wire _al_u1654_o;
  wire _al_u1656_o;
  wire _al_u1657_o;
  wire _al_u1658_o;
  wire _al_u1659_o;
  wire _al_u1660_o;
  wire _al_u1662_o;
  wire _al_u1663_o;
  wire _al_u1664_o;
  wire _al_u1667_o;
  wire _al_u1668_o;
  wire _al_u1670_o;
  wire _al_u1675_o;
  wire _al_u1676_o;
  wire _al_u1679_o;
  wire _al_u1681_o;
  wire _al_u1683_o;
  wire _al_u1685_o;
  wire _al_u1687_o;
  wire _al_u1689_o;
  wire _al_u1690_o;
  wire _al_u1692_o;
  wire _al_u1694_o;
  wire _al_u1695_o;
  wire _al_u1697_o;
  wire _al_u1699_o;
  wire _al_u1701_o;
  wire _al_u1703_o;
  wire _al_u1704_o;
  wire _al_u1706_o;
  wire _al_u1708_o;
  wire _al_u1710_o;
  wire _al_u1712_o;
  wire _al_u1713_o;
  wire _al_u1715_o;
  wire _al_u1716_o;
  wire _al_u1718_o;
  wire _al_u1720_o;
  wire _al_u1721_o;
  wire _al_u1723_o;
  wire _al_u1724_o;
  wire _al_u1726_o;
  wire _al_u1727_o;
  wire _al_u1730_o;
  wire _al_u1733_o;
  wire _al_u1734_o;
  wire _al_u1737_o;
  wire _al_u1741_o;
  wire _al_u1743_o;
  wire _al_u1749_o;
  wire _al_u1751_o;
  wire _al_u1752_o;
  wire _al_u1753_o;
  wire _al_u1755_o;
  wire _al_u1756_o;
  wire _al_u1757_o;
  wire _al_u1758_o;
  wire _al_u1759_o;
  wire _al_u1761_o;
  wire _al_u1762_o;
  wire _al_u1763_o;
  wire _al_u1765_o;
  wire _al_u1767_o;
  wire _al_u1768_o;
  wire _al_u1769_o;
  wire _al_u1770_o;
  wire _al_u1772_o;
  wire _al_u1774_o;
  wire _al_u1775_o;
  wire _al_u1777_o;
  wire _al_u1778_o;
  wire _al_u1779_o;
  wire _al_u1781_o;
  wire _al_u1782_o;
  wire _al_u1783_o;
  wire _al_u1784_o;
  wire _al_u1785_o;
  wire _al_u1787_o;
  wire _al_u1788_o;
  wire _al_u1791_o;
  wire _al_u1793_o;
  wire _al_u1794_o;
  wire _al_u1796_o;
  wire _al_u1797_o;
  wire _al_u1799_o;
  wire _al_u1801_o;
  wire _al_u1802_o;
  wire _al_u1803_o;
  wire _al_u1804_o;
  wire _al_u1806_o;
  wire _al_u1808_o;
  wire _al_u1809_o;
  wire _al_u1810_o;
  wire _al_u1811_o;
  wire _al_u1812_o;
  wire _al_u1813_o;
  wire _al_u1815_o;
  wire _al_u1816_o;
  wire _al_u1817_o;
  wire _al_u1818_o;
  wire _al_u1819_o;
  wire _al_u1820_o;
  wire _al_u1821_o;
  wire _al_u1823_o;
  wire _al_u1824_o;
  wire _al_u1826_o;
  wire _al_u1827_o;
  wire _al_u1829_o;
  wire _al_u1830_o;
  wire _al_u1832_o;
  wire _al_u1833_o;
  wire _al_u1835_o;
  wire _al_u1836_o;
  wire _al_u1838_o;
  wire _al_u1839_o;
  wire _al_u1841_o;
  wire _al_u1843_o;
  wire _al_u1844_o;
  wire _al_u1846_o;
  wire _al_u1848_o;
  wire _al_u1850_o;
  wire _al_u1852_o;
  wire _al_u1854_o;
  wire _al_u1856_o;
  wire _al_u1858_o;
  wire _al_u1859_o;
  wire _al_u1861_o;
  wire _al_u1862_o;
  wire _al_u1864_o;
  wire _al_u1865_o;
  wire _al_u1867_o;
  wire _al_u1868_o;
  wire _al_u1875_o;
  wire _al_u1881_o;
  wire _al_u1882_o;
  wire _al_u1883_o;
  wire _al_u1885_o;
  wire _al_u1886_o;
  wire _al_u1887_o;
  wire _al_u1888_o;
  wire _al_u1891_o;
  wire _al_u1892_o;
  wire _al_u1893_o;
  wire _al_u1894_o;
  wire _al_u1895_o;
  wire _al_u1896_o;
  wire _al_u1899_o;
  wire _al_u1900_o;
  wire _al_u1902_o;
  wire _al_u1905_o;
  wire _al_u1906_o;
  wire _al_u1907_o;
  wire _al_u1910_o;
  wire _al_u1911_o;
  wire _al_u1912_o;
  wire _al_u1913_o;
  wire _al_u1915_o;
  wire _al_u1916_o;
  wire _al_u1917_o;
  wire _al_u1919_o;
  wire _al_u1920_o;
  wire _al_u1921_o;
  wire _al_u1923_o;
  wire _al_u1924_o;
  wire _al_u1925_o;
  wire _al_u1926_o;
  wire _al_u1928_o;
  wire _al_u1929_o;
  wire _al_u1930_o;
  wire _al_u1932_o;
  wire _al_u1933_o;
  wire _al_u1934_o;
  wire _al_u1935_o;
  wire _al_u1937_o;
  wire _al_u1938_o;
  wire _al_u1939_o;
  wire _al_u1941_o;
  wire _al_u1942_o;
  wire _al_u1943_o;
  wire _al_u1944_o;
  wire _al_u1946_o;
  wire _al_u1947_o;
  wire _al_u1948_o;
  wire _al_u1950_o;
  wire _al_u1951_o;
  wire _al_u1952_o;
  wire _al_u1953_o;
  wire _al_u1955_o;
  wire _al_u1956_o;
  wire _al_u1957_o;
  wire _al_u1959_o;
  wire _al_u1960_o;
  wire _al_u1961_o;
  wire _al_u1962_o;
  wire _al_u1964_o;
  wire _al_u1965_o;
  wire _al_u1966_o;
  wire _al_u1967_o;
  wire _al_u1968_o;
  wire _al_u1969_o;
  wire _al_u1971_o;
  wire _al_u1972_o;
  wire _al_u1973_o;
  wire _al_u1974_o;
  wire _al_u1975_o;
  wire _al_u1976_o;
  wire _al_u1977_o;
  wire _al_u1979_o;
  wire _al_u1982_o;
  wire _al_u1983_o;
  wire _al_u1986_o;
  wire _al_u1987_o;
  wire _al_u1988_o;
  wire _al_u1993_o;
  wire _al_u2032_o;
  wire _al_u2033_o;
  wire _al_u2034_o;
  wire _al_u2035_o;
  wire _al_u2036_o;
  wire _al_u2037_o;
  wire _al_u2038_o;
  wire _al_u2040_o;
  wire _al_u2055_o;
  wire _al_u2056_o;
  wire _al_u2057_o;
  wire _al_u2059_o;
  wire _al_u2060_o;
  wire _al_u2061_o;
  wire _al_u2062_o;
  wire _al_u2063_o;
  wire _al_u2077_o;
  wire _al_u2078_o;
  wire _al_u2079_o;
  wire _al_u2080_o;
  wire _al_u2081_o;
  wire _al_u2082_o;
  wire _al_u2083_o;
  wire _al_u2084_o;
  wire _al_u2085_o;
  wire _al_u2099_o;
  wire _al_u2100_o;
  wire _al_u2101_o;
  wire _al_u2102_o;
  wire _al_u2104_o;
  wire _al_u2105_o;
  wire _al_u2106_o;
  wire _al_u2107_o;
  wire _al_u2121_o;
  wire _al_u2122_o;
  wire _al_u2123_o;
  wire _al_u2124_o;
  wire _al_u2125_o;
  wire _al_u2126_o;
  wire _al_u2127_o;
  wire _al_u2128_o;
  wire _al_u2129_o;
  wire _al_u2143_o;
  wire _al_u2144_o;
  wire _al_u2145_o;
  wire _al_u2146_o;
  wire _al_u2148_o;
  wire _al_u2149_o;
  wire _al_u2150_o;
  wire _al_u2151_o;
  wire _al_u2165_o;
  wire _al_u2166_o;
  wire _al_u2167_o;
  wire _al_u2168_o;
  wire _al_u2170_o;
  wire _al_u2171_o;
  wire _al_u2173_o;
  wire _al_u2201_o;
  wire _al_u2202_o;
  wire _al_u2203_o;
  wire _al_u2204_o;
  wire _al_u2205_o;
  wire _al_u2207_o;
  wire _al_u2208_o;
  wire _al_u2210_o;
  wire _al_u2211_o;
  wire _al_u2212_o;
  wire _al_u2213_o;
  wire _al_u2215_o;
  wire _al_u2216_o;
  wire _al_u2217_o;
  wire _al_u2219_o;
  wire _al_u2220_o;
  wire _al_u2221_o;
  wire _al_u2223_o;
  wire _al_u2224_o;
  wire _al_u2225_o;
  wire _al_u2228_o;
  wire _al_u2229_o;
  wire _al_u2230_o;
  wire _al_u2231_o;
  wire _al_u2233_o;
  wire _al_u2234_o;
  wire _al_u2235_o;
  wire _al_u2237_o;
  wire _al_u2238_o;
  wire _al_u2239_o;
  wire _al_u2240_o;
  wire _al_u2242_o;
  wire _al_u2243_o;
  wire _al_u2244_o;
  wire _al_u2246_o;
  wire _al_u2247_o;
  wire _al_u2248_o;
  wire _al_u2250_o;
  wire _al_u2251_o;
  wire _al_u2252_o;
  wire _al_u2255_o;
  wire _al_u2256_o;
  wire _al_u2257_o;
  wire _al_u2259_o;
  wire _al_u2260_o;
  wire _al_u2261_o;
  wire _al_u2262_o;
  wire _al_u2264_o;
  wire _al_u2265_o;
  wire _al_u2266_o;
  wire _al_u2267_o;
  wire _al_u2268_o;
  wire _al_u2269_o;
  wire _al_u2270_o;
  wire _al_u2272_o;
  wire _al_u2274_o;
  wire _al_u2275_o;
  wire _al_u2276_o;
  wire _al_u2277_o;
  wire _al_u2278_o;
  wire _al_u2279_o;
  wire _al_u2280_o;
  wire _al_u2281_o;
  wire _al_u2283_o;
  wire _al_u2284_o;
  wire _al_u2285_o;
  wire _al_u2288_o;
  wire _al_u2289_o;
  wire _al_u2290_o;
  wire _al_u2292_o;
  wire _al_u2293_o;
  wire _al_u2295_o;
  wire _al_u2296_o;
  wire _al_u2297_o;
  wire _al_u2298_o;
  wire _al_u2299_o;
  wire _al_u2305_o;
  wire _al_u2306_o;
  wire _al_u2309_o;
  wire _al_u2312_o;
  wire _al_u2315_o;
  wire _al_u2317_o;
  wire _al_u2319_o;
  wire _al_u2321_o;
  wire _al_u2323_o;
  wire _al_u2325_o;
  wire _al_u2327_o;
  wire _al_u2329_o;
  wire _al_u2331_o;
  wire _al_u2333_o;
  wire _al_u2335_o;
  wire _al_u2337_o;
  wire _al_u2339_o;
  wire _al_u2341_o;
  wire _al_u2343_o;
  wire _al_u2345_o;
  wire _al_u2347_o;
  wire _al_u2349_o;
  wire _al_u2351_o;
  wire _al_u2353_o;
  wire _al_u2355_o;
  wire _al_u2357_o;
  wire _al_u2359_o;
  wire _al_u2361_o;
  wire _al_u2364_o;
  wire _al_u2365_o;
  wire _al_u2366_o;
  wire _al_u2367_o;
  wire _al_u2369_o;
  wire _al_u2370_o;
  wire _al_u2371_o;
  wire _al_u2373_o;
  wire _al_u2375_o;
  wire _al_u2376_o;
  wire _al_u2377_o;
  wire _al_u2378_o;
  wire _al_u2379_o;
  wire _al_u2380_o;
  wire _al_u2381_o;
  wire _al_u2382_o;
  wire _al_u2386_o;
  wire _al_u2387_o;
  wire _al_u2388_o;
  wire _al_u2389_o;
  wire _al_u2390_o;
  wire _al_u2392_o;
  wire _al_u2393_o;
  wire _al_u2395_o;
  wire _al_u2396_o;
  wire _al_u2397_o;
  wire _al_u2398_o;
  wire _al_u2399_o;
  wire _al_u2403_o;
  wire _al_u2404_o;
  wire _al_u2405_o;
  wire _al_u2406_o;
  wire _al_u2407_o;
  wire _al_u2409_o;
  wire _al_u2411_o;
  wire _al_u2412_o;
  wire _al_u2413_o;
  wire _al_u2414_o;
  wire _al_u2415_o;
  wire _al_u2416_o;
  wire _al_u2417_o;
  wire _al_u2418_o;
  wire _al_u2419_o;
  wire _al_u2420_o;
  wire _al_u2423_o;
  wire _al_u2424_o;
  wire _al_u2425_o;
  wire _al_u2426_o;
  wire _al_u2427_o;
  wire _al_u2428_o;
  wire _al_u2429_o;
  wire _al_u2433_o;
  wire _al_u2434_o;
  wire _al_u2435_o;
  wire _al_u2437_o;
  wire _al_u2438_o;
  wire _al_u2439_o;
  wire _al_u2441_o;
  wire _al_u2442_o;
  wire _al_u2443_o;
  wire _al_u2445_o;
  wire _al_u2446_o;
  wire _al_u2447_o;
  wire _al_u2449_o;
  wire _al_u2450_o;
  wire _al_u2451_o;
  wire _al_u2453_o;
  wire _al_u2454_o;
  wire _al_u2455_o;
  wire _al_u2458_o;
  wire _al_u2459_o;
  wire _al_u2460_o;
  wire _al_u2461_o;
  wire _al_u2463_o;
  wire _al_u2464_o;
  wire _al_u2467_o;
  wire _al_u2468_o;
  wire _al_u2469_o;
  wire _al_u2470_o;
  wire _al_u2476_o;
  wire _al_u2478_o;
  wire _al_u2480_o;
  wire _al_u2482_o;
  wire _al_u2484_o;
  wire _al_u2488_o;
  wire _al_u2490_o;
  wire _al_u2492_o;
  wire _al_u2494_o;
  wire _al_u2496_o;
  wire _al_u2500_o;
  wire _al_u2502_o;
  wire _al_u2504_o;
  wire _al_u2506_o;
  wire _al_u2508_o;
  wire _al_u2512_o;
  wire _al_u2514_o;
  wire _al_u2516_o;
  wire _al_u2518_o;
  wire _al_u2520_o;
  wire _al_u2642_o;
  wire _al_u2643_o;
  wire _al_u2644_o;
  wire _al_u2646_o;
  wire _al_u2647_o;
  wire _al_u2648_o;
  wire _al_u2649_o;
  wire _al_u2650_o;
  wire _al_u2717_o;
  wire _al_u2721_o;
  wire _al_u2724_o;
  wire _al_u2725_o;
  wire _al_u2728_o;
  wire _al_u2729_o;
  wire _al_u2733_o;
  wire _al_u2740_o;
  wire _al_u2741_o;
  wire _al_u2746_o;
  wire _al_u2747_o;
  wire _al_u2748_o;
  wire _al_u2749_o;
  wire _al_u2750_o;
  wire _al_u2751_o;
  wire _al_u2754_o;
  wire _al_u2755_o;
  wire _al_u2756_o;
  wire _al_u2758_o;
  wire _al_u2759_o;
  wire _al_u2760_o;
  wire _al_u2761_o;
  wire _al_u2763_o;
  wire _al_u2764_o;
  wire _al_u2766_o;
  wire _al_u2767_o;
  wire _al_u2770_o;
  wire _al_u2771_o;
  wire _al_u2772_o;
  wire _al_u2773_o;
  wire _al_u2774_o;
  wire _al_u2776_o;
  wire _al_u2778_o;
  wire _al_u2779_o;
  wire _al_u2782_o;
  wire _al_u2783_o;
  wire _al_u2784_o;
  wire _al_u2785_o;
  wire _al_u2786_o;
  wire _al_u2787_o;
  wire _al_u2789_o;
  wire _al_u2790_o;
  wire _al_u2791_o;
  wire _al_u2793_o;
  wire _al_u2794_o;
  wire _al_u2800_o;
  wire _al_u2802_o;
  wire _al_u2803_o;
  wire _al_u2804_o;
  wire _al_u2808_o;
  wire _al_u2809_o;
  wire _al_u2810_o;
  wire _al_u2813_o;
  wire _al_u2815_o;
  wire _al_u2816_o;
  wire _al_u2817_o;
  wire _al_u2818_o;
  wire _al_u2824_o;
  wire _al_u2825_o;
  wire _al_u2827_o;
  wire _al_u2829_o;
  wire _al_u2832_o;
  wire _al_u2834_o;
  wire _al_u2835_o;
  wire _al_u2836_o;
  wire _al_u2837_o;
  wire _al_u2839_o;
  wire _al_u2840_o;
  wire _al_u2841_o;
  wire _al_u2843_o;
  wire _al_u2845_o;
  wire _al_u2846_o;
  wire _al_u2847_o;
  wire _al_u2849_o;
  wire _al_u2855_o;
  wire _al_u2857_o;
  wire _al_u2858_o;
  wire _al_u2860_o;
  wire _al_u2861_o;
  wire _al_u2862_o;
  wire _al_u2863_o;
  wire _al_u2865_o;
  wire _al_u2866_o;
  wire _al_u2867_o;
  wire _al_u2868_o;
  wire _al_u2869_o;
  wire _al_u2870_o;
  wire _al_u2871_o;
  wire _al_u2872_o;
  wire _al_u2873_o;
  wire _al_u2875_o;
  wire _al_u2877_o;
  wire _al_u2878_o;
  wire _al_u2881_o;
  wire _al_u2882_o;
  wire _al_u2920_o;
  wire _al_u2921_o;
  wire _al_u2937_o;
  wire _al_u2953_o;
  wire _al_u2969_o;
  wire _al_u2985_o;
  wire _al_u2986_o;
  wire _al_u2988_o;
  wire _al_u2990_o;
  wire _al_u2992_o;
  wire _al_u3000_o;
  wire _al_u3002_o;
  wire _al_u3004_o;
  wire _al_u3006_o;
  wire _al_u3008_o;
  wire _al_u3010_o;
  wire _al_u3012_o;
  wire _al_u3015_o;
  wire _al_u3017_o;
  wire _al_u3020_o;
  wire _al_u3021_o;
  wire _al_u3022_o;
  wire _al_u3023_o;
  wire _al_u3024_o;
  wire _al_u3026_o;
  wire _al_u3027_o;
  wire _al_u3029_o;
  wire _al_u3030_o;
  wire _al_u3032_o;
  wire _al_u3034_o;
  wire _al_u3035_o;
  wire _al_u3040_o;
  wire _al_u3041_o;
  wire _al_u3046_o;
  wire _al_u3047_o;
  wire _al_u3052_o;
  wire _al_u3053_o;
  wire _al_u3057_o;
  wire _al_u3058_o;
  wire _al_u3062_o;
  wire _al_u3063_o;
  wire _al_u3067_o;
  wire _al_u3068_o;
  wire _al_u3072_o;
  wire _al_u3073_o;
  wire _al_u3075_o;
  wire _al_u3076_o;
  wire _al_u3078_o;
  wire _al_u3079_o;
  wire _al_u3080_o;
  wire _al_u3081_o;
  wire _al_u3082_o;
  wire _al_u3083_o;
  wire _al_u3085_o;
  wire _al_u3086_o;
  wire _al_u3087_o;
  wire _al_u3091_o;
  wire _al_u3092_o;
  wire _al_u3094_o;
  wire _al_u3096_o;
  wire _al_u3097_o;
  wire _al_u3100_o;
  wire _al_u3101_o;
  wire _al_u3102_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3105_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3108_o;
  wire _al_u3109_o;
  wire _al_u3110_o;
  wire _al_u3111_o;
  wire _al_u3114_o;
  wire _al_u3115_o;
  wire _al_u3117_o;
  wire _al_u3118_o;
  wire _al_u3119_o;
  wire _al_u3120_o;
  wire _al_u3121_o;
  wire _al_u3122_o;
  wire _al_u3124_o;
  wire _al_u3126_o;
  wire _al_u3127_o;
  wire _al_u3129_o;
  wire _al_u3132_o;
  wire _al_u3133_o;
  wire _al_u3148_o;
  wire _al_u3149_o;
  wire _al_u3150_o;
  wire _al_u3151_o;
  wire _al_u3152_o;
  wire _al_u3156_o;
  wire _al_u3157_o;
  wire _al_u3158_o;
  wire _al_u3159_o;
  wire _al_u3160_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3166_o;
  wire _al_u3167_o;
  wire _al_u3169_o;
  wire _al_u3170_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3175_o;
  wire _al_u3176_o;
  wire _al_u3179_o;
  wire _al_u3180_o;
  wire _al_u3181_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3193_o;
  wire _al_u3196_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3199_o;
  wire _al_u3201_o;
  wire _al_u3202_o;
  wire _al_u3203_o;
  wire _al_u3205_o;
  wire _al_u3206_o;
  wire _al_u3208_o;
  wire _al_u3210_o;
  wire _al_u3211_o;
  wire _al_u3214_o;
  wire _al_u3215_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3218_o;
  wire _al_u3219_o;
  wire _al_u3221_o;
  wire _al_u3222_o;
  wire _al_u3223_o;
  wire _al_u3224_o;
  wire _al_u3225_o;
  wire _al_u3226_o;
  wire _al_u3227_o;
  wire _al_u3229_o;
  wire _al_u3230_o;
  wire _al_u3233_o;
  wire _al_u3234_o;
  wire _al_u3235_o;
  wire _al_u3236_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3239_o;
  wire _al_u3240_o;
  wire _al_u3242_o;
  wire _al_u3243_o;
  wire _al_u3245_o;
  wire _al_u3246_o;
  wire _al_u3248_o;
  wire _al_u3249_o;
  wire _al_u3255_o;
  wire _al_u3256_o;
  wire _al_u3258_o;
  wire _al_u3259_o;
  wire _al_u3268_o;
  wire _al_u3270_o;
  wire _al_u3271_o;
  wire _al_u3274_o;
  wire _al_u3275_o;
  wire _al_u3279_o;
  wire _al_u3280_o;
  wire _al_u3281_o;
  wire _al_u3286_o;
  wire _al_u3287_o;
  wire _al_u3305_o;
  wire _al_u3306_o;
  wire _al_u3307_o;
  wire _al_u3308_o;
  wire _al_u3309_o;
  wire _al_u3312_o;
  wire _al_u3313_o;
  wire _al_u3314_o;
  wire _al_u3318_o;
  wire _al_u3319_o;
  wire _al_u3320_o;
  wire _al_u3322_o;
  wire _al_u3323_o;
  wire _al_u3324_o;
  wire _al_u3325_o;
  wire _al_u3326_o;
  wire _al_u3327_o;
  wire _al_u3328_o;
  wire _al_u3329_o;
  wire _al_u3333_o;
  wire _al_u3334_o;
  wire _al_u3335_o;
  wire _al_u3337_o;
  wire _al_u3338_o;
  wire _al_u3339_o;
  wire _al_u3342_o;
  wire _al_u3343_o;
  wire _al_u3345_o;
  wire _al_u3348_o;
  wire _al_u3350_o;
  wire _al_u3352_o;
  wire _al_u3355_o;
  wire _al_u3356_o;
  wire _al_u3357_o;
  wire _al_u3358_o;
  wire _al_u3359_o;
  wire _al_u3360_o;
  wire _al_u3361_o;
  wire _al_u3365_o;
  wire _al_u3366_o;
  wire _al_u3367_o;
  wire _al_u3368_o;
  wire _al_u3369_o;
  wire _al_u3370_o;
  wire _al_u3371_o;
  wire _al_u3372_o;
  wire _al_u3378_o;
  wire _al_u3381_o;
  wire _al_u3384_o;
  wire _al_u3385_o;
  wire _al_u3387_o;
  wire _al_u3388_o;
  wire _al_u3390_o;
  wire _al_u3391_o;
  wire _al_u3392_o;
  wire _al_u3393_o;
  wire _al_u3395_o;
  wire _al_u3396_o;
  wire _al_u3397_o;
  wire _al_u3398_o;
  wire _al_u3399_o;
  wire _al_u3400_o;
  wire _al_u3401_o;
  wire _al_u3402_o;
  wire _al_u3405_o;
  wire _al_u3410_o;
  wire _al_u3414_o;
  wire _al_u3415_o;
  wire _al_u3416_o;
  wire _al_u3419_o;
  wire _al_u3420_o;
  wire _al_u3421_o;
  wire _al_u3422_o;
  wire _al_u3423_o;
  wire _al_u3424_o;
  wire _al_u3429_o;
  wire _al_u3430_o;
  wire _al_u3431_o;
  wire _al_u3434_o;
  wire _al_u3435_o;
  wire _al_u3438_o;
  wire _al_u3439_o;
  wire _al_u3440_o;
  wire _al_u3441_o;
  wire _al_u3442_o;
  wire _al_u3443_o;
  wire _al_u3445_o;
  wire _al_u3446_o;
  wire _al_u3448_o;
  wire _al_u3449_o;
  wire _al_u3450_o;
  wire _al_u3451_o;
  wire _al_u3453_o;
  wire _al_u3454_o;
  wire _al_u3456_o;
  wire _al_u3457_o;
  wire _al_u3460_o;
  wire _al_u3461_o;
  wire _al_u3462_o;
  wire _al_u3463_o;
  wire _al_u3465_o;
  wire _al_u3466_o;
  wire _al_u3467_o;
  wire _al_u3468_o;
  wire _al_u3470_o;
  wire _al_u3471_o;
  wire _al_u3472_o;
  wire _al_u3473_o;
  wire _al_u3476_o;
  wire _al_u3477_o;
  wire _al_u3478_o;
  wire _al_u3479_o;
  wire _al_u3481_o;
  wire _al_u3482_o;
  wire _al_u3483_o;
  wire _al_u3486_o;
  wire _al_u3487_o;
  wire _al_u3488_o;
  wire _al_u3489_o;
  wire _al_u3491_o;
  wire _al_u3492_o;
  wire _al_u3493_o;
  wire _al_u3494_o;
  wire _al_u3497_o;
  wire _al_u3498_o;
  wire _al_u3499_o;
  wire _al_u3502_o;
  wire _al_u3503_o;
  wire _al_u3504_o;
  wire _al_u3507_o;
  wire _al_u3508_o;
  wire _al_u3509_o;
  wire _al_u3512_o;
  wire _al_u3513_o;
  wire _al_u3514_o;
  wire _al_u3515_o;
  wire _al_u3517_o;
  wire _al_u3518_o;
  wire _al_u3519_o;
  wire _al_u3520_o;
  wire _al_u3522_o;
  wire _al_u3523_o;
  wire _al_u3524_o;
  wire _al_u3527_o;
  wire _al_u3528_o;
  wire _al_u3529_o;
  wire _al_u3530_o;
  wire _al_u3532_o;
  wire _al_u3533_o;
  wire _al_u3534_o;
  wire _al_u3535_o;
  wire _al_u3538_o;
  wire _al_u3539_o;
  wire _al_u3540_o;
  wire _al_u3542_o;
  wire _al_u3544_o;
  wire _al_u3547_o;
  wire _al_u3549_o;
  wire _al_u3552_o;
  wire _al_u3553_o;
  wire _al_u3554_o;
  wire _al_u3555_o;
  wire _al_u3556_o;
  wire _al_u3557_o;
  wire _al_u3558_o;
  wire _al_u3559_o;
  wire _al_u355_o;
  wire _al_u3560_o;
  wire _al_u3561_o;
  wire _al_u3562_o;
  wire _al_u3563_o;
  wire _al_u3564_o;
  wire _al_u3565_o;
  wire _al_u3568_o;
  wire _al_u3569_o;
  wire _al_u3570_o;
  wire _al_u3571_o;
  wire _al_u3573_o;
  wire _al_u3574_o;
  wire _al_u3575_o;
  wire _al_u3576_o;
  wire _al_u3578_o;
  wire _al_u3579_o;
  wire _al_u357_o;
  wire _al_u3580_o;
  wire _al_u3581_o;
  wire _al_u3582_o;
  wire _al_u3583_o;
  wire _al_u3584_o;
  wire _al_u3585_o;
  wire _al_u3586_o;
  wire _al_u3587_o;
  wire _al_u3588_o;
  wire _al_u358_o;
  wire _al_u3591_o;
  wire _al_u3592_o;
  wire _al_u3593_o;
  wire _al_u3596_o;
  wire _al_u3597_o;
  wire _al_u359_o;
  wire _al_u3601_o;
  wire _al_u3603_o;
  wire _al_u3608_o;
  wire _al_u3609_o;
  wire _al_u360_o;
  wire _al_u3610_o;
  wire _al_u3611_o;
  wire _al_u3612_o;
  wire _al_u3613_o;
  wire _al_u3614_o;
  wire _al_u3615_o;
  wire _al_u3617_o;
  wire _al_u3618_o;
  wire _al_u3620_o;
  wire _al_u3621_o;
  wire _al_u3622_o;
  wire _al_u3624_o;
  wire _al_u3625_o;
  wire _al_u3626_o;
  wire _al_u3627_o;
  wire _al_u3628_o;
  wire _al_u3629_o;
  wire _al_u3630_o;
  wire _al_u3631_o;
  wire _al_u3632_o;
  wire _al_u3633_o;
  wire _al_u3634_o;
  wire _al_u3635_o;
  wire _al_u3636_o;
  wire _al_u3637_o;
  wire _al_u3638_o;
  wire _al_u3639_o;
  wire _al_u3640_o;
  wire _al_u3641_o;
  wire _al_u3643_o;
  wire _al_u3646_o;
  wire _al_u3647_o;
  wire _al_u3648_o;
  wire _al_u3649_o;
  wire _al_u364_o;
  wire _al_u3650_o;
  wire _al_u3652_o;
  wire _al_u3653_o;
  wire _al_u3654_o;
  wire _al_u3655_o;
  wire _al_u3657_o;
  wire _al_u3658_o;
  wire _al_u3659_o;
  wire _al_u3661_o;
  wire _al_u3662_o;
  wire _al_u3663_o;
  wire _al_u3664_o;
  wire _al_u3665_o;
  wire _al_u3666_o;
  wire _al_u3667_o;
  wire _al_u3669_o;
  wire _al_u3670_o;
  wire _al_u3672_o;
  wire _al_u3673_o;
  wire _al_u3674_o;
  wire _al_u3675_o;
  wire _al_u3677_o;
  wire _al_u3678_o;
  wire _al_u3679_o;
  wire _al_u367_o;
  wire _al_u3680_o;
  wire _al_u3681_o;
  wire _al_u3683_o;
  wire _al_u3684_o;
  wire _al_u3686_o;
  wire _al_u3688_o;
  wire _al_u368_o;
  wire _al_u3690_o;
  wire _al_u3691_o;
  wire _al_u3692_o;
  wire _al_u3693_o;
  wire _al_u3694_o;
  wire _al_u3695_o;
  wire _al_u3696_o;
  wire _al_u3697_o;
  wire _al_u3699_o;
  wire _al_u3700_o;
  wire _al_u3701_o;
  wire _al_u3702_o;
  wire _al_u3703_o;
  wire _al_u3704_o;
  wire _al_u3705_o;
  wire _al_u3706_o;
  wire _al_u3707_o;
  wire _al_u3708_o;
  wire _al_u3709_o;
  wire _al_u370_o;
  wire _al_u3710_o;
  wire _al_u3713_o;
  wire _al_u3715_o;
  wire _al_u3716_o;
  wire _al_u3717_o;
  wire _al_u3718_o;
  wire _al_u3719_o;
  wire _al_u3720_o;
  wire _al_u3721_o;
  wire _al_u3722_o;
  wire _al_u3724_o;
  wire _al_u3725_o;
  wire _al_u3726_o;
  wire _al_u3727_o;
  wire _al_u3728_o;
  wire _al_u3729_o;
  wire _al_u3730_o;
  wire _al_u3731_o;
  wire _al_u3732_o;
  wire _al_u3733_o;
  wire _al_u3734_o;
  wire _al_u3735_o;
  wire _al_u3736_o;
  wire _al_u3738_o;
  wire _al_u3739_o;
  wire _al_u3740_o;
  wire _al_u3741_o;
  wire _al_u3742_o;
  wire _al_u3743_o;
  wire _al_u3744_o;
  wire _al_u3745_o;
  wire _al_u3747_o;
  wire _al_u3748_o;
  wire _al_u3749_o;
  wire _al_u374_o;
  wire _al_u3750_o;
  wire _al_u3753_o;
  wire _al_u3754_o;
  wire _al_u3755_o;
  wire _al_u3758_o;
  wire _al_u3769_o;
  wire _al_u3776_o;
  wire _al_u3777_o;
  wire _al_u3779_o;
  wire _al_u3780_o;
  wire _al_u3781_o;
  wire _al_u3782_o;
  wire _al_u3783_o;
  wire _al_u3784_o;
  wire _al_u3787_o;
  wire _al_u3788_o;
  wire _al_u3789_o;
  wire _al_u3790_o;
  wire _al_u3791_o;
  wire _al_u3792_o;
  wire _al_u3793_o;
  wire _al_u3794_o;
  wire _al_u3795_o;
  wire _al_u3796_o;
  wire _al_u3797_o;
  wire _al_u3798_o;
  wire _al_u3799_o;
  wire _al_u379_o;
  wire _al_u3800_o;
  wire _al_u3801_o;
  wire _al_u3803_o;
  wire _al_u3804_o;
  wire _al_u3805_o;
  wire _al_u3806_o;
  wire _al_u3807_o;
  wire _al_u3808_o;
  wire _al_u3810_o;
  wire _al_u3811_o;
  wire _al_u3812_o;
  wire _al_u3813_o;
  wire _al_u3814_o;
  wire _al_u3815_o;
  wire _al_u3816_o;
  wire _al_u3817_o;
  wire _al_u3818_o;
  wire _al_u3819_o;
  wire _al_u3820_o;
  wire _al_u3821_o;
  wire _al_u3822_o;
  wire _al_u3823_o;
  wire _al_u3824_o;
  wire _al_u3825_o;
  wire _al_u3826_o;
  wire _al_u3827_o;
  wire _al_u3829_o;
  wire _al_u3830_o;
  wire _al_u3831_o;
  wire _al_u3832_o;
  wire _al_u3833_o;
  wire _al_u3834_o;
  wire _al_u3835_o;
  wire _al_u3836_o;
  wire _al_u3837_o;
  wire _al_u3838_o;
  wire _al_u3839_o;
  wire _al_u3840_o;
  wire _al_u3841_o;
  wire _al_u3843_o;
  wire _al_u3844_o;
  wire _al_u3845_o;
  wire _al_u3846_o;
  wire _al_u3847_o;
  wire _al_u3848_o;
  wire _al_u3849_o;
  wire _al_u3851_o;
  wire _al_u3853_o;
  wire _al_u3854_o;
  wire _al_u3855_o;
  wire _al_u3856_o;
  wire _al_u3857_o;
  wire _al_u3858_o;
  wire _al_u3859_o;
  wire _al_u3869_o;
  wire _al_u3870_o;
  wire _al_u3872_o;
  wire _al_u3874_o;
  wire _al_u3875_o;
  wire _al_u3878_o;
  wire _al_u3879_o;
  wire _al_u3880_o;
  wire _al_u3882_o;
  wire _al_u3884_o;
  wire _al_u3885_o;
  wire _al_u3887_o;
  wire _al_u3889_o;
  wire _al_u388_o;
  wire _al_u3891_o;
  wire _al_u3892_o;
  wire _al_u3893_o;
  wire _al_u3894_o;
  wire _al_u3895_o;
  wire _al_u3896_o;
  wire _al_u3897_o;
  wire _al_u3898_o;
  wire _al_u3900_o;
  wire _al_u3901_o;
  wire _al_u3902_o;
  wire _al_u3903_o;
  wire _al_u3904_o;
  wire _al_u3905_o;
  wire _al_u3906_o;
  wire _al_u3907_o;
  wire _al_u3908_o;
  wire _al_u3909_o;
  wire _al_u3910_o;
  wire _al_u3911_o;
  wire _al_u3912_o;
  wire _al_u3914_o;
  wire _al_u3915_o;
  wire _al_u3916_o;
  wire _al_u3917_o;
  wire _al_u3918_o;
  wire _al_u3919_o;
  wire _al_u3920_o;
  wire _al_u3921_o;
  wire _al_u3922_o;
  wire _al_u3924_o;
  wire _al_u3925_o;
  wire _al_u3926_o;
  wire _al_u3927_o;
  wire _al_u3929_o;
  wire _al_u3931_o;
  wire _al_u3932_o;
  wire _al_u3934_o;
  wire _al_u3935_o;
  wire _al_u3937_o;
  wire _al_u3938_o;
  wire _al_u3940_o;
  wire _al_u3941_o;
  wire _al_u3943_o;
  wire _al_u3944_o;
  wire _al_u3946_o;
  wire _al_u3947_o;
  wire _al_u3949_o;
  wire _al_u3950_o;
  wire _al_u3952_o;
  wire _al_u3953_o;
  wire _al_u3955_o;
  wire _al_u3956_o;
  wire _al_u3958_o;
  wire _al_u3959_o;
  wire _al_u3961_o;
  wire _al_u3962_o;
  wire _al_u3964_o;
  wire _al_u3966_o;
  wire _al_u3967_o;
  wire _al_u3969_o;
  wire _al_u3970_o;
  wire _al_u3972_o;
  wire _al_u3973_o;
  wire _al_u3975_o;
  wire _al_u3976_o;
  wire _al_u3978_o;
  wire _al_u3979_o;
  wire _al_u3981_o;
  wire _al_u3982_o;
  wire _al_u3984_o;
  wire _al_u3985_o;
  wire _al_u3987_o;
  wire _al_u3988_o;
  wire _al_u3990_o;
  wire _al_u3991_o;
  wire _al_u3993_o;
  wire _al_u3994_o;
  wire _al_u3995_o;
  wire _al_u3996_o;
  wire _al_u3997_o;
  wire _al_u4000_o;
  wire _al_u4001_o;
  wire _al_u4002_o;
  wire _al_u4003_o;
  wire _al_u4004_o;
  wire _al_u4007_o;
  wire _al_u4008_o;
  wire _al_u4009_o;
  wire _al_u4010_o;
  wire _al_u4011_o;
  wire _al_u4012_o;
  wire _al_u4013_o;
  wire _al_u4014_o;
  wire _al_u4015_o;
  wire _al_u4016_o;
  wire _al_u4017_o;
  wire _al_u4018_o;
  wire _al_u4019_o;
  wire _al_u4021_o;
  wire _al_u4022_o;
  wire _al_u4023_o;
  wire _al_u4025_o;
  wire _al_u4027_o;
  wire _al_u4028_o;
  wire _al_u4029_o;
  wire _al_u4030_o;
  wire _al_u4031_o;
  wire _al_u4032_o;
  wire _al_u4034_o;
  wire _al_u4035_o;
  wire _al_u4036_o;
  wire _al_u4037_o;
  wire _al_u4038_o;
  wire _al_u4039_o;
  wire _al_u4040_o;
  wire _al_u4041_o;
  wire _al_u4042_o;
  wire _al_u4043_o;
  wire _al_u4044_o;
  wire _al_u4045_o;
  wire _al_u4046_o;
  wire _al_u4048_o;
  wire _al_u4049_o;
  wire _al_u4052_o;
  wire _al_u4055_o;
  wire _al_u4056_o;
  wire _al_u4058_o;
  wire _al_u405_o;
  wire _al_u4060_o;
  wire _al_u4061_o;
  wire _al_u4063_o;
  wire _al_u4065_o;
  wire _al_u4066_o;
  wire _al_u4068_o;
  wire _al_u4070_o;
  wire _al_u4071_o;
  wire _al_u4073_o;
  wire _al_u4075_o;
  wire _al_u4076_o;
  wire _al_u4078_o;
  wire _al_u4080_o;
  wire _al_u4081_o;
  wire _al_u4083_o;
  wire _al_u4085_o;
  wire _al_u4086_o;
  wire _al_u4088_o;
  wire _al_u4090_o;
  wire _al_u4091_o;
  wire _al_u4093_o;
  wire _al_u4095_o;
  wire _al_u4096_o;
  wire _al_u4098_o;
  wire _al_u4100_o;
  wire _al_u4101_o;
  wire _al_u4103_o;
  wire _al_u4105_o;
  wire _al_u4106_o;
  wire _al_u4108_o;
  wire _al_u4110_o;
  wire _al_u4111_o;
  wire _al_u4113_o;
  wire _al_u4115_o;
  wire _al_u4116_o;
  wire _al_u4118_o;
  wire _al_u4120_o;
  wire _al_u4121_o;
  wire _al_u4123_o;
  wire _al_u4125_o;
  wire _al_u4126_o;
  wire _al_u4128_o;
  wire _al_u4130_o;
  wire _al_u4131_o;
  wire _al_u4133_o;
  wire _al_u4135_o;
  wire _al_u4136_o;
  wire _al_u4138_o;
  wire _al_u4140_o;
  wire _al_u4141_o;
  wire _al_u4143_o;
  wire _al_u4145_o;
  wire _al_u4146_o;
  wire _al_u4147_o;
  wire _al_u4148_o;
  wire _al_u4150_o;
  wire _al_u4151_o;
  wire _al_u4152_o;
  wire _al_u4153_o;
  wire _al_u4154_o;
  wire _al_u4155_o;
  wire _al_u4156_o;
  wire _al_u4157_o;
  wire _al_u4158_o;
  wire _al_u4159_o;
  wire _al_u4160_o;
  wire _al_u4161_o;
  wire _al_u4162_o;
  wire _al_u4163_o;
  wire _al_u4164_o;
  wire _al_u4165_o;
  wire _al_u4166_o;
  wire _al_u4168_o;
  wire _al_u4169_o;
  wire _al_u4170_o;
  wire _al_u4171_o;
  wire _al_u4172_o;
  wire _al_u4173_o;
  wire _al_u4175_o;
  wire _al_u4181_o;
  wire _al_u4182_o;
  wire _al_u4183_o;
  wire _al_u4184_o;
  wire _al_u4188_o;
  wire _al_u4189_o;
  wire _al_u4190_o;
  wire _al_u4191_o;
  wire _al_u4194_o;
  wire _al_u4195_o;
  wire _al_u4196_o;
  wire _al_u4197_o;
  wire _al_u4200_o;
  wire _al_u4201_o;
  wire _al_u4204_o;
  wire _al_u4205_o;
  wire _al_u4208_o;
  wire _al_u4209_o;
  wire _al_u4212_o;
  wire _al_u4213_o;
  wire _al_u4216_o;
  wire _al_u4217_o;
  wire _al_u4218_o;
  wire _al_u4219_o;
  wire _al_u4222_o;
  wire _al_u4223_o;
  wire _al_u4224_o;
  wire _al_u4225_o;
  wire _al_u4228_o;
  wire _al_u4229_o;
  wire _al_u4230_o;
  wire _al_u4231_o;
  wire _al_u4234_o;
  wire _al_u4235_o;
  wire _al_u4236_o;
  wire _al_u4237_o;
  wire _al_u4239_o;
  wire _al_u4240_o;
  wire _al_u4242_o;
  wire _al_u4243_o;
  wire _al_u4244_o;
  wire _al_u4245_o;
  wire _al_u4246_o;
  wire _al_u4247_o;
  wire _al_u4248_o;
  wire _al_u4249_o;
  wire _al_u4251_o;
  wire _al_u4252_o;
  wire _al_u4256_o;
  wire _al_u4258_o;
  wire _al_u4259_o;
  wire _al_u4260_o;
  wire _al_u4261_o;
  wire _al_u4262_o;
  wire _al_u4263_o;
  wire _al_u4266_o;
  wire _al_u4267_o;
  wire _al_u4269_o;
  wire _al_u4271_o;
  wire _al_u4272_o;
  wire _al_u4273_o;
  wire _al_u4274_o;
  wire _al_u4278_o;
  wire _al_u4280_o;
  wire _al_u4281_o;
  wire _al_u4282_o;
  wire _al_u4283_o;
  wire _al_u4284_o;
  wire _al_u4289_o;
  wire _al_u4290_o;
  wire _al_u4291_o;
  wire _al_u4292_o;
  wire _al_u4293_o;
  wire _al_u4294_o;
  wire _al_u4295_o;
  wire _al_u4297_o;
  wire _al_u4300_o;
  wire _al_u4302_o;
  wire _al_u4304_o;
  wire _al_u4305_o;
  wire _al_u4306_o;
  wire _al_u4308_o;
  wire _al_u4309_o;
  wire _al_u4310_o;
  wire _al_u4311_o;
  wire _al_u4312_o;
  wire _al_u4313_o;
  wire _al_u4314_o;
  wire _al_u4315_o;
  wire _al_u4316_o;
  wire _al_u4317_o;
  wire _al_u4318_o;
  wire _al_u4319_o;
  wire _al_u4320_o;
  wire _al_u4322_o;
  wire _al_u4323_o;
  wire _al_u4324_o;
  wire _al_u4325_o;
  wire _al_u4326_o;
  wire _al_u4327_o;
  wire _al_u4328_o;
  wire _al_u4329_o;
  wire _al_u4330_o;
  wire _al_u4331_o;
  wire _al_u4332_o;
  wire _al_u4333_o;
  wire _al_u4334_o;
  wire _al_u4336_o;
  wire _al_u4337_o;
  wire _al_u4338_o;
  wire _al_u4339_o;
  wire _al_u4340_o;
  wire _al_u4341_o;
  wire _al_u4342_o;
  wire _al_u4343_o;
  wire _al_u4344_o;
  wire _al_u4345_o;
  wire _al_u4346_o;
  wire _al_u4350_o;
  wire _al_u4351_o;
  wire _al_u4352_o;
  wire _al_u4353_o;
  wire _al_u4354_o;
  wire _al_u4355_o;
  wire _al_u4356_o;
  wire _al_u4357_o;
  wire _al_u4358_o;
  wire _al_u4359_o;
  wire _al_u4360_o;
  wire _al_u4361_o;
  wire _al_u4362_o;
  wire _al_u4363_o;
  wire _al_u4364_o;
  wire _al_u4367_o;
  wire _al_u4368_o;
  wire _al_u4371_o;
  wire _al_u4372_o;
  wire _al_u4373_o;
  wire _al_u4374_o;
  wire _al_u4375_o;
  wire _al_u4376_o;
  wire _al_u4377_o;
  wire _al_u4378_o;
  wire _al_u4379_o;
  wire _al_u4380_o;
  wire _al_u4381_o;
  wire _al_u4382_o;
  wire _al_u4383_o;
  wire _al_u4384_o;
  wire _al_u4385_o;
  wire _al_u4386_o;
  wire _al_u4387_o;
  wire _al_u4388_o;
  wire _al_u4389_o;
  wire _al_u4390_o;
  wire _al_u4391_o;
  wire _al_u4392_o;
  wire _al_u4393_o;
  wire _al_u4395_o;
  wire _al_u4396_o;
  wire _al_u4397_o;
  wire _al_u4398_o;
  wire _al_u4399_o;
  wire _al_u4400_o;
  wire _al_u4401_o;
  wire _al_u4402_o;
  wire _al_u4403_o;
  wire _al_u4404_o;
  wire _al_u4405_o;
  wire _al_u4406_o;
  wire _al_u4407_o;
  wire _al_u4408_o;
  wire _al_u4409_o;
  wire _al_u4410_o;
  wire _al_u4411_o;
  wire _al_u4412_o;
  wire _al_u4413_o;
  wire _al_u4414_o;
  wire _al_u4415_o;
  wire _al_u4416_o;
  wire _al_u4419_o;
  wire _al_u4421_o;
  wire _al_u4422_o;
  wire _al_u4423_o;
  wire _al_u4425_o;
  wire _al_u4426_o;
  wire _al_u4438_o;
  wire _al_u4450_o;
  wire _al_u4451_o;
  wire _al_u4452_o;
  wire _al_u4455_o;
  wire _al_u4456_o;
  wire _al_u4457_o;
  wire _al_u4459_o;
  wire _al_u4460_o;
  wire _al_u4461_o;
  wire _al_u4462_o;
  wire _al_u4463_o;
  wire _al_u4464_o;
  wire _al_u4465_o;
  wire _al_u4466_o;
  wire _al_u4467_o;
  wire _al_u4468_o;
  wire _al_u4470_o;
  wire _al_u4471_o;
  wire _al_u4472_o;
  wire _al_u4473_o;
  wire _al_u4474_o;
  wire _al_u4475_o;
  wire _al_u4476_o;
  wire _al_u4478_o;
  wire _al_u4480_o;
  wire _al_u4481_o;
  wire _al_u4483_o;
  wire _al_u4484_o;
  wire _al_u4485_o;
  wire _al_u4486_o;
  wire _al_u4487_o;
  wire _al_u4488_o;
  wire _al_u4490_o;
  wire _al_u4492_o;
  wire _al_u4495_o;
  wire _al_u4499_o;
  wire _al_u4500_o;
  wire _al_u4501_o;
  wire _al_u4509_o;
  wire _al_u4511_o;
  wire _al_u4512_o;
  wire _al_u4513_o;
  wire _al_u4514_o;
  wire _al_u4515_o;
  wire _al_u4516_o;
  wire _al_u4517_o;
  wire _al_u4519_o;
  wire _al_u4520_o;
  wire _al_u4521_o;
  wire _al_u4523_o;
  wire _al_u4524_o;
  wire _al_u4525_o;
  wire _al_u4526_o;
  wire _al_u4527_o;
  wire _al_u4528_o;
  wire _al_u4529_o;
  wire _al_u452_o;
  wire _al_u4530_o;
  wire _al_u4532_o;
  wire _al_u4533_o;
  wire _al_u4534_o;
  wire _al_u4535_o;
  wire _al_u4537_o;
  wire _al_u4539_o;
  wire _al_u453_o;
  wire _al_u4542_o;
  wire _al_u4544_o;
  wire _al_u4545_o;
  wire _al_u4546_o;
  wire _al_u4548_o;
  wire _al_u4549_o;
  wire _al_u4550_o;
  wire _al_u4551_o;
  wire _al_u4552_o;
  wire _al_u4553_o;
  wire _al_u4557_o;
  wire _al_u4558_o;
  wire _al_u4559_o;
  wire _al_u4560_o;
  wire _al_u4561_o;
  wire _al_u4562_o;
  wire _al_u4563_o;
  wire _al_u4564_o;
  wire _al_u4566_o;
  wire _al_u4567_o;
  wire _al_u4568_o;
  wire _al_u4569_o;
  wire _al_u456_o;
  wire _al_u4571_o;
  wire _al_u4573_o;
  wire _al_u4574_o;
  wire _al_u4575_o;
  wire _al_u4576_o;
  wire _al_u4577_o;
  wire _al_u4578_o;
  wire _al_u4580_o;
  wire _al_u4581_o;
  wire _al_u4582_o;
  wire _al_u4583_o;
  wire _al_u4584_o;
  wire _al_u4586_o;
  wire _al_u4587_o;
  wire _al_u4588_o;
  wire _al_u4589_o;
  wire _al_u4591_o;
  wire _al_u4592_o;
  wire _al_u4593_o;
  wire _al_u4594_o;
  wire _al_u4595_o;
  wire _al_u4596_o;
  wire _al_u4597_o;
  wire _al_u4598_o;
  wire _al_u4599_o;
  wire _al_u4600_o;
  wire _al_u4601_o;
  wire _al_u4602_o;
  wire _al_u4603_o;
  wire _al_u4604_o;
  wire _al_u4605_o;
  wire _al_u4607_o;
  wire _al_u4608_o;
  wire _al_u4609_o;
  wire _al_u4610_o;
  wire _al_u4611_o;
  wire _al_u4612_o;
  wire _al_u4613_o;
  wire _al_u4616_o;
  wire _al_u4617_o;
  wire _al_u4618_o;
  wire _al_u4619_o;
  wire _al_u4620_o;
  wire _al_u4621_o;
  wire _al_u4623_o;
  wire _al_u4624_o;
  wire _al_u4625_o;
  wire _al_u4626_o;
  wire _al_u4627_o;
  wire _al_u4628_o;
  wire _al_u4629_o;
  wire _al_u462_o;
  wire _al_u4631_o;
  wire _al_u4633_o;
  wire _al_u4634_o;
  wire _al_u4635_o;
  wire _al_u4636_o;
  wire _al_u4637_o;
  wire _al_u4638_o;
  wire _al_u4639_o;
  wire _al_u463_o;
  wire _al_u4642_o;
  wire _al_u4643_o;
  wire _al_u4644_o;
  wire _al_u4645_o;
  wire _al_u4646_o;
  wire _al_u4647_o;
  wire _al_u4649_o;
  wire _al_u4650_o;
  wire _al_u4651_o;
  wire _al_u4652_o;
  wire _al_u4653_o;
  wire _al_u4654_o;
  wire _al_u4655_o;
  wire _al_u4657_o;
  wire _al_u4659_o;
  wire _al_u465_o;
  wire _al_u4660_o;
  wire _al_u4661_o;
  wire _al_u4662_o;
  wire _al_u4663_o;
  wire _al_u4664_o;
  wire _al_u4665_o;
  wire _al_u4668_o;
  wire _al_u4669_o;
  wire _al_u4670_o;
  wire _al_u4671_o;
  wire _al_u4672_o;
  wire _al_u4673_o;
  wire _al_u4675_o;
  wire _al_u4676_o;
  wire _al_u4677_o;
  wire _al_u4678_o;
  wire _al_u4679_o;
  wire _al_u467_o;
  wire _al_u4680_o;
  wire _al_u4681_o;
  wire _al_u4682_o;
  wire _al_u4683_o;
  wire _al_u4684_o;
  wire _al_u4685_o;
  wire _al_u4686_o;
  wire _al_u4687_o;
  wire _al_u4688_o;
  wire _al_u4689_o;
  wire _al_u4690_o;
  wire _al_u4692_o;
  wire _al_u4693_o;
  wire _al_u4694_o;
  wire _al_u4695_o;
  wire _al_u4697_o;
  wire _al_u4698_o;
  wire _al_u4699_o;
  wire _al_u4700_o;
  wire _al_u4701_o;
  wire _al_u4702_o;
  wire _al_u4703_o;
  wire _al_u4704_o;
  wire _al_u4705_o;
  wire _al_u4706_o;
  wire _al_u4708_o;
  wire _al_u4709_o;
  wire _al_u470_o;
  wire _al_u4711_o;
  wire _al_u4712_o;
  wire _al_u4713_o;
  wire _al_u4716_o;
  wire _al_u4717_o;
  wire _al_u4718_o;
  wire _al_u4719_o;
  wire _al_u4720_o;
  wire _al_u4722_o;
  wire _al_u4723_o;
  wire _al_u4724_o;
  wire _al_u4725_o;
  wire _al_u4726_o;
  wire _al_u4727_o;
  wire _al_u4728_o;
  wire _al_u4729_o;
  wire _al_u472_o;
  wire _al_u4730_o;
  wire _al_u4731_o;
  wire _al_u4732_o;
  wire _al_u4733_o;
  wire _al_u4734_o;
  wire _al_u4735_o;
  wire _al_u4736_o;
  wire _al_u4737_o;
  wire _al_u473_o;
  wire _al_u4740_o;
  wire _al_u4741_o;
  wire _al_u4742_o;
  wire _al_u4743_o;
  wire _al_u4744_o;
  wire _al_u4746_o;
  wire _al_u4747_o;
  wire _al_u4749_o;
  wire _al_u4750_o;
  wire _al_u4751_o;
  wire _al_u4752_o;
  wire _al_u4753_o;
  wire _al_u4754_o;
  wire _al_u4755_o;
  wire _al_u4756_o;
  wire _al_u4757_o;
  wire _al_u4758_o;
  wire _al_u475_o;
  wire _al_u4760_o;
  wire _al_u4761_o;
  wire _al_u4762_o;
  wire _al_u4763_o;
  wire _al_u4764_o;
  wire _al_u4766_o;
  wire _al_u4767_o;
  wire _al_u4768_o;
  wire _al_u4769_o;
  wire _al_u4770_o;
  wire _al_u4772_o;
  wire _al_u4773_o;
  wire _al_u4774_o;
  wire _al_u4775_o;
  wire _al_u4776_o;
  wire _al_u4777_o;
  wire _al_u4780_o;
  wire _al_u4781_o;
  wire _al_u4782_o;
  wire _al_u4783_o;
  wire _al_u4784_o;
  wire _al_u4786_o;
  wire _al_u4787_o;
  wire _al_u4788_o;
  wire _al_u4789_o;
  wire _al_u478_o;
  wire _al_u4790_o;
  wire _al_u4792_o;
  wire _al_u4793_o;
  wire _al_u4794_o;
  wire _al_u4795_o;
  wire _al_u4796_o;
  wire _al_u4797_o;
  wire _al_u4801_o;
  wire _al_u4802_o;
  wire _al_u4803_o;
  wire _al_u4804_o;
  wire _al_u4805_o;
  wire _al_u4806_o;
  wire _al_u4807_o;
  wire _al_u4808_o;
  wire _al_u4809_o;
  wire _al_u480_o;
  wire _al_u4810_o;
  wire _al_u4811_o;
  wire _al_u4812_o;
  wire _al_u4814_o;
  wire _al_u4815_o;
  wire _al_u4816_o;
  wire _al_u4817_o;
  wire _al_u481_o;
  wire _al_u4820_o;
  wire _al_u4821_o;
  wire _al_u4822_o;
  wire _al_u4823_o;
  wire _al_u4824_o;
  wire _al_u4826_o;
  wire _al_u4827_o;
  wire _al_u4828_o;
  wire _al_u4829_o;
  wire _al_u482_o;
  wire _al_u4830_o;
  wire _al_u4832_o;
  wire _al_u4833_o;
  wire _al_u4834_o;
  wire _al_u4835_o;
  wire _al_u4836_o;
  wire _al_u4837_o;
  wire _al_u4838_o;
  wire _al_u483_o;
  wire _al_u4841_o;
  wire _al_u4842_o;
  wire _al_u4844_o;
  wire _al_u4845_o;
  wire _al_u4846_o;
  wire _al_u4847_o;
  wire _al_u4848_o;
  wire _al_u4849_o;
  wire _al_u4850_o;
  wire _al_u4851_o;
  wire _al_u4852_o;
  wire _al_u4853_o;
  wire _al_u4854_o;
  wire _al_u4855_o;
  wire _al_u4857_o;
  wire _al_u4858_o;
  wire _al_u4859_o;
  wire _al_u4860_o;
  wire _al_u4861_o;
  wire _al_u4862_o;
  wire _al_u4863_o;
  wire _al_u4865_o;
  wire _al_u4866_o;
  wire _al_u4867_o;
  wire _al_u486_o;
  wire _al_u4871_o;
  wire _al_u4872_o;
  wire _al_u4873_o;
  wire _al_u4874_o;
  wire _al_u4875_o;
  wire _al_u4876_o;
  wire _al_u4877_o;
  wire _al_u4878_o;
  wire _al_u4879_o;
  wire _al_u487_o;
  wire _al_u4880_o;
  wire _al_u4881_o;
  wire _al_u4882_o;
  wire _al_u4884_o;
  wire _al_u4885_o;
  wire _al_u4886_o;
  wire _al_u4887_o;
  wire _al_u488_o;
  wire _al_u4890_o;
  wire _al_u4891_o;
  wire _al_u4892_o;
  wire _al_u4893_o;
  wire _al_u4894_o;
  wire _al_u4896_o;
  wire _al_u4897_o;
  wire _al_u4898_o;
  wire _al_u489_o;
  wire _al_u4900_o;
  wire _al_u4901_o;
  wire _al_u4902_o;
  wire _al_u4903_o;
  wire _al_u4904_o;
  wire _al_u4905_o;
  wire _al_u4906_o;
  wire _al_u4908_o;
  wire _al_u4909_o;
  wire _al_u4910_o;
  wire _al_u4912_o;
  wire _al_u4914_o;
  wire _al_u4916_o;
  wire _al_u4917_o;
  wire _al_u4918_o;
  wire _al_u4919_o;
  wire _al_u491_o;
  wire _al_u4920_o;
  wire _al_u4921_o;
  wire _al_u4922_o;
  wire _al_u4923_o;
  wire _al_u4925_o;
  wire _al_u4927_o;
  wire _al_u4928_o;
  wire _al_u492_o;
  wire _al_u4930_o;
  wire _al_u4931_o;
  wire _al_u4932_o;
  wire _al_u4934_o;
  wire _al_u4935_o;
  wire _al_u4937_o;
  wire _al_u4938_o;
  wire _al_u4939_o;
  wire _al_u493_o;
  wire _al_u4940_o;
  wire _al_u4941_o;
  wire _al_u4942_o;
  wire _al_u4943_o;
  wire _al_u4944_o;
  wire _al_u4945_o;
  wire _al_u4946_o;
  wire _al_u4947_o;
  wire _al_u4948_o;
  wire _al_u4949_o;
  wire _al_u494_o;
  wire _al_u4950_o;
  wire _al_u4951_o;
  wire _al_u4953_o;
  wire _al_u4954_o;
  wire _al_u4955_o;
  wire _al_u4957_o;
  wire _al_u4959_o;
  wire _al_u4961_o;
  wire _al_u4963_o;
  wire _al_u4965_o;
  wire _al_u4967_o;
  wire _al_u4969_o;
  wire _al_u496_o;
  wire _al_u4970_o;
  wire _al_u4971_o;
  wire _al_u4973_o;
  wire _al_u4974_o;
  wire _al_u4975_o;
  wire _al_u4977_o;
  wire _al_u497_o;
  wire _al_u4981_o;
  wire _al_u4982_o;
  wire _al_u4983_o;
  wire _al_u4984_o;
  wire _al_u4985_o;
  wire _al_u4986_o;
  wire _al_u4987_o;
  wire _al_u4988_o;
  wire _al_u4989_o;
  wire _al_u498_o;
  wire _al_u4990_o;
  wire _al_u4993_o;
  wire _al_u4994_o;
  wire _al_u499_o;
  wire _al_u5000_o;
  wire _al_u5001_o;
  wire _al_u5003_o;
  wire _al_u5006_o;
  wire _al_u5009_o;
  wire _al_u5017_o;
  wire _al_u5020_o;
  wire _al_u5021_o;
  wire _al_u5023_o;
  wire _al_u5024_o;
  wire _al_u5025_o;
  wire _al_u5026_o;
  wire _al_u5028_o;
  wire _al_u5029_o;
  wire _al_u5030_o;
  wire _al_u5031_o;
  wire _al_u5032_o;
  wire _al_u5036_o;
  wire _al_u5037_o;
  wire _al_u5038_o;
  wire _al_u5039_o;
  wire _al_u5040_o;
  wire _al_u5044_o;
  wire _al_u5047_o;
  wire _al_u5048_o;
  wire _al_u5049_o;
  wire _al_u5050_o;
  wire _al_u5051_o;
  wire _al_u5052_o;
  wire _al_u5053_o;
  wire _al_u5055_o;
  wire _al_u5056_o;
  wire _al_u5057_o;
  wire _al_u5058_o;
  wire _al_u5059_o;
  wire _al_u5061_o;
  wire _al_u5062_o;
  wire _al_u5063_o;
  wire _al_u5066_o;
  wire _al_u5067_o;
  wire _al_u5069_o;
  wire _al_u5070_o;
  wire _al_u5071_o;
  wire _al_u5072_o;
  wire _al_u5073_o;
  wire _al_u5074_o;
  wire _al_u5075_o;
  wire _al_u5076_o;
  wire _al_u5078_o;
  wire _al_u5080_o;
  wire _al_u5081_o;
  wire _al_u5082_o;
  wire _al_u5083_o;
  wire _al_u5084_o;
  wire _al_u5085_o;
  wire _al_u5086_o;
  wire _al_u5087_o;
  wire _al_u5088_o;
  wire _al_u5090_o;
  wire _al_u5091_o;
  wire _al_u5092_o;
  wire _al_u5094_o;
  wire _al_u5095_o;
  wire _al_u5096_o;
  wire _al_u5097_o;
  wire _al_u5098_o;
  wire _al_u5099_o;
  wire _al_u5100_o;
  wire _al_u5101_o;
  wire _al_u5103_o;
  wire _al_u5104_o;
  wire _al_u5105_o;
  wire _al_u5107_o;
  wire _al_u5108_o;
  wire _al_u5109_o;
  wire _al_u5110_o;
  wire _al_u5111_o;
  wire _al_u5112_o;
  wire _al_u5113_o;
  wire _al_u5114_o;
  wire _al_u5116_o;
  wire _al_u5117_o;
  wire _al_u5118_o;
  wire _al_u5119_o;
  wire _al_u5120_o;
  wire _al_u5121_o;
  wire _al_u5122_o;
  wire _al_u5125_o;
  wire _al_u5126_o;
  wire _al_u5127_o;
  wire _al_u5128_o;
  wire _al_u5130_o;
  wire _al_u5131_o;
  wire _al_u5132_o;
  wire _al_u5133_o;
  wire _al_u5134_o;
  wire _al_u5135_o;
  wire _al_u5136_o;
  wire _al_u5137_o;
  wire _al_u5138_o;
  wire _al_u5139_o;
  wire _al_u5140_o;
  wire _al_u5141_o;
  wire _al_u5142_o;
  wire _al_u5143_o;
  wire _al_u5144_o;
  wire _al_u5145_o;
  wire _al_u5146_o;
  wire _al_u5147_o;
  wire _al_u5148_o;
  wire _al_u5149_o;
  wire _al_u5151_o;
  wire _al_u5152_o;
  wire _al_u5153_o;
  wire _al_u5154_o;
  wire _al_u5156_o;
  wire _al_u5157_o;
  wire _al_u5159_o;
  wire _al_u5163_o;
  wire _al_u5164_o;
  wire _al_u5165_o;
  wire _al_u5166_o;
  wire _al_u5167_o;
  wire _al_u5168_o;
  wire _al_u5169_o;
  wire _al_u5171_o;
  wire _al_u5173_o;
  wire _al_u5176_o;
  wire _al_u5177_o;
  wire _al_u5178_o;
  wire _al_u5179_o;
  wire _al_u5180_o;
  wire _al_u5181_o;
  wire _al_u5183_o;
  wire _al_u5186_o;
  wire _al_u5187_o;
  wire _al_u5188_o;
  wire _al_u5189_o;
  wire _al_u5190_o;
  wire _al_u5191_o;
  wire _al_u5192_o;
  wire _al_u5193_o;
  wire _al_u5194_o;
  wire _al_u5196_o;
  wire _al_u5197_o;
  wire _al_u5198_o;
  wire _al_u5199_o;
  wire _al_u5200_o;
  wire _al_u5201_o;
  wire _al_u5203_o;
  wire _al_u5204_o;
  wire _al_u5206_o;
  wire _al_u5207_o;
  wire _al_u5208_o;
  wire _al_u5213_o;
  wire _al_u5214_o;
  wire _al_u5215_o;
  wire _al_u5216_o;
  wire _al_u5217_o;
  wire _al_u5218_o;
  wire _al_u5219_o;
  wire _al_u5220_o;
  wire _al_u5222_o;
  wire _al_u5223_o;
  wire _al_u5224_o;
  wire _al_u5225_o;
  wire _al_u5229_o;
  wire _al_u5230_o;
  wire _al_u5231_o;
  wire _al_u5232_o;
  wire _al_u5233_o;
  wire _al_u5235_o;
  wire _al_u5236_o;
  wire _al_u5237_o;
  wire _al_u5238_o;
  wire _al_u5239_o;
  wire _al_u5240_o;
  wire _al_u5241_o;
  wire _al_u5242_o;
  wire _al_u5243_o;
  wire _al_u5245_o;
  wire _al_u5246_o;
  wire _al_u5251_o;
  wire _al_u5252_o;
  wire _al_u5253_o;
  wire _al_u5254_o;
  wire _al_u5255_o;
  wire _al_u5256_o;
  wire _al_u5257_o;
  wire _al_u5258_o;
  wire _al_u5260_o;
  wire _al_u5261_o;
  wire _al_u5262_o;
  wire _al_u5263_o;
  wire _al_u5264_o;
  wire _al_u5265_o;
  wire _al_u5266_o;
  wire _al_u5267_o;
  wire _al_u5268_o;
  wire _al_u526_o;
  wire _al_u5271_o;
  wire _al_u5274_o;
  wire _al_u5275_o;
  wire _al_u5276_o;
  wire _al_u5278_o;
  wire _al_u5280_o;
  wire _al_u5282_o;
  wire _al_u5284_o;
  wire _al_u5285_o;
  wire _al_u5286_o;
  wire _al_u5287_o;
  wire _al_u5288_o;
  wire _al_u5291_o;
  wire _al_u5292_o;
  wire _al_u5293_o;
  wire _al_u5294_o;
  wire _al_u5295_o;
  wire _al_u5296_o;
  wire _al_u5297_o;
  wire _al_u5298_o;
  wire _al_u5299_o;
  wire _al_u529_o;
  wire _al_u5300_o;
  wire _al_u5301_o;
  wire _al_u5302_o;
  wire _al_u5303_o;
  wire _al_u5304_o;
  wire _al_u5305_o;
  wire _al_u5307_o;
  wire _al_u5308_o;
  wire _al_u530_o;
  wire _al_u5310_o;
  wire _al_u5311_o;
  wire _al_u5312_o;
  wire _al_u5313_o;
  wire _al_u5315_o;
  wire _al_u5316_o;
  wire _al_u5317_o;
  wire _al_u5318_o;
  wire _al_u5319_o;
  wire _al_u5320_o;
  wire _al_u5321_o;
  wire _al_u5323_o;
  wire _al_u5324_o;
  wire _al_u5325_o;
  wire _al_u5327_o;
  wire _al_u5328_o;
  wire _al_u5329_o;
  wire _al_u5331_o;
  wire _al_u5332_o;
  wire _al_u5333_o;
  wire _al_u5334_o;
  wire _al_u5335_o;
  wire _al_u5336_o;
  wire _al_u5337_o;
  wire _al_u5338_o;
  wire _al_u5339_o;
  wire _al_u533_o;
  wire _al_u5340_o;
  wire _al_u5341_o;
  wire _al_u5344_o;
  wire _al_u5345_o;
  wire _al_u5346_o;
  wire _al_u5347_o;
  wire _al_u5348_o;
  wire _al_u5349_o;
  wire _al_u5351_o;
  wire _al_u5352_o;
  wire _al_u5353_o;
  wire _al_u5354_o;
  wire _al_u5355_o;
  wire _al_u5357_o;
  wire _al_u5358_o;
  wire _al_u5359_o;
  wire _al_u5360_o;
  wire _al_u5361_o;
  wire _al_u5362_o;
  wire _al_u5364_o;
  wire _al_u5365_o;
  wire _al_u5366_o;
  wire _al_u5369_o;
  wire _al_u5370_o;
  wire _al_u5371_o;
  wire _al_u5375_o;
  wire _al_u5376_o;
  wire _al_u5377_o;
  wire _al_u5378_o;
  wire _al_u5379_o;
  wire _al_u5380_o;
  wire _al_u5381_o;
  wire _al_u5382_o;
  wire _al_u5383_o;
  wire _al_u5384_o;
  wire _al_u5385_o;
  wire _al_u5386_o;
  wire _al_u5387_o;
  wire _al_u5389_o;
  wire _al_u5390_o;
  wire _al_u5392_o;
  wire _al_u5394_o;
  wire _al_u5395_o;
  wire _al_u5396_o;
  wire _al_u5398_o;
  wire _al_u5399_o;
  wire _al_u5400_o;
  wire _al_u5403_o;
  wire _al_u5407_o;
  wire _al_u5408_o;
  wire _al_u540_o;
  wire _al_u5411_o;
  wire _al_u5412_o;
  wire _al_u5413_o;
  wire _al_u5415_o;
  wire _al_u5416_o;
  wire _al_u5417_o;
  wire _al_u5419_o;
  wire _al_u5420_o;
  wire _al_u5421_o;
  wire _al_u5424_o;
  wire _al_u5425_o;
  wire _al_u5426_o;
  wire _al_u5428_o;
  wire _al_u5429_o;
  wire _al_u5430_o;
  wire _al_u5431_o;
  wire _al_u5433_o;
  wire _al_u5435_o;
  wire _al_u5437_o;
  wire _al_u5438_o;
  wire _al_u5439_o;
  wire _al_u543_o;
  wire _al_u5441_o;
  wire _al_u5442_o;
  wire _al_u5444_o;
  wire _al_u5445_o;
  wire _al_u5446_o;
  wire _al_u5448_o;
  wire _al_u5449_o;
  wire _al_u544_o;
  wire _al_u5451_o;
  wire _al_u5452_o;
  wire _al_u5453_o;
  wire _al_u5454_o;
  wire _al_u5455_o;
  wire _al_u5457_o;
  wire _al_u5458_o;
  wire _al_u5460_o;
  wire _al_u5462_o;
  wire _al_u5463_o;
  wire _al_u5465_o;
  wire _al_u5466_o;
  wire _al_u5467_o;
  wire _al_u5468_o;
  wire _al_u546_o;
  wire _al_u5470_o;
  wire _al_u5471_o;
  wire _al_u5473_o;
  wire _al_u5474_o;
  wire _al_u5476_o;
  wire _al_u5477_o;
  wire _al_u5478_o;
  wire _al_u5479_o;
  wire _al_u5481_o;
  wire _al_u5482_o;
  wire _al_u5484_o;
  wire _al_u5485_o;
  wire _al_u5486_o;
  wire _al_u5487_o;
  wire _al_u5488_o;
  wire _al_u5489_o;
  wire _al_u5493_o;
  wire _al_u5495_o;
  wire _al_u5497_o;
  wire _al_u5498_o;
  wire _al_u5499_o;
  wire _al_u5501_o;
  wire _al_u5504_o;
  wire _al_u5505_o;
  wire _al_u5507_o;
  wire _al_u5508_o;
  wire _al_u5510_o;
  wire _al_u5511_o;
  wire _al_u5513_o;
  wire _al_u5514_o;
  wire _al_u5515_o;
  wire _al_u5516_o;
  wire _al_u5518_o;
  wire _al_u5519_o;
  wire _al_u5520_o;
  wire _al_u5522_o;
  wire _al_u5523_o;
  wire _al_u5524_o;
  wire _al_u552_o;
  wire _al_u5531_o;
  wire _al_u5532_o;
  wire _al_u5533_o;
  wire _al_u5534_o;
  wire _al_u5536_o;
  wire _al_u5537_o;
  wire _al_u5539_o;
  wire _al_u553_o;
  wire _al_u5541_o;
  wire _al_u5542_o;
  wire _al_u5544_o;
  wire _al_u5546_o;
  wire _al_u5547_o;
  wire _al_u5549_o;
  wire _al_u554_o;
  wire _al_u5550_o;
  wire _al_u5552_o;
  wire _al_u5553_o;
  wire _al_u5554_o;
  wire _al_u5556_o;
  wire _al_u5558_o;
  wire _al_u5559_o;
  wire _al_u555_o;
  wire _al_u5561_o;
  wire _al_u5562_o;
  wire _al_u5564_o;
  wire _al_u5565_o;
  wire _al_u5567_o;
  wire _al_u5568_o;
  wire _al_u556_o;
  wire _al_u5570_o;
  wire _al_u5571_o;
  wire _al_u5573_o;
  wire _al_u5574_o;
  wire _al_u5575_o;
  wire _al_u5577_o;
  wire _al_u5578_o;
  wire _al_u557_o;
  wire _al_u5580_o;
  wire _al_u5581_o;
  wire _al_u5582_o;
  wire _al_u5583_o;
  wire _al_u5584_o;
  wire _al_u5585_o;
  wire _al_u5587_o;
  wire _al_u5588_o;
  wire _al_u5590_o;
  wire _al_u5591_o;
  wire _al_u5592_o;
  wire _al_u5593_o;
  wire _al_u5594_o;
  wire _al_u5595_o;
  wire _al_u5597_o;
  wire _al_u5598_o;
  wire _al_u5599_o;
  wire _al_u5600_o;
  wire _al_u5601_o;
  wire _al_u5603_o;
  wire _al_u5604_o;
  wire _al_u5605_o;
  wire _al_u5607_o;
  wire _al_u5608_o;
  wire _al_u5609_o;
  wire _al_u560_o;
  wire _al_u5614_o;
  wire _al_u5616_o;
  wire _al_u5618_o;
  wire _al_u5619_o;
  wire _al_u5620_o;
  wire _al_u5622_o;
  wire _al_u5623_o;
  wire _al_u5625_o;
  wire _al_u5626_o;
  wire _al_u5629_o;
  wire _al_u5632_o;
  wire _al_u5633_o;
  wire _al_u5635_o;
  wire _al_u5636_o;
  wire _al_u5637_o;
  wire _al_u5638_o;
  wire _al_u5643_o;
  wire _al_u5644_o;
  wire _al_u5647_o;
  wire _al_u5648_o;
  wire _al_u5649_o;
  wire _al_u5650_o;
  wire _al_u5651_o;
  wire _al_u5652_o;
  wire _al_u5654_o;
  wire _al_u5655_o;
  wire _al_u5656_o;
  wire _al_u5657_o;
  wire _al_u5658_o;
  wire _al_u5659_o;
  wire _al_u5660_o;
  wire _al_u5661_o;
  wire _al_u5663_o;
  wire _al_u5664_o;
  wire _al_u5665_o;
  wire _al_u5666_o;
  wire _al_u5667_o;
  wire _al_u5668_o;
  wire _al_u566_o;
  wire _al_u5670_o;
  wire _al_u5671_o;
  wire _al_u5672_o;
  wire _al_u5673_o;
  wire _al_u5674_o;
  wire _al_u5675_o;
  wire _al_u5676_o;
  wire _al_u5677_o;
  wire _al_u5678_o;
  wire _al_u5679_o;
  wire _al_u5680_o;
  wire _al_u5682_o;
  wire _al_u5683_o;
  wire _al_u5684_o;
  wire _al_u5685_o;
  wire _al_u5687_o;
  wire _al_u5688_o;
  wire _al_u5689_o;
  wire _al_u5690_o;
  wire _al_u5692_o;
  wire _al_u5693_o;
  wire _al_u5694_o;
  wire _al_u5695_o;
  wire _al_u5696_o;
  wire _al_u5697_o;
  wire _al_u5698_o;
  wire _al_u5699_o;
  wire _al_u569_o;
  wire _al_u5700_o;
  wire _al_u5701_o;
  wire _al_u5702_o;
  wire _al_u5704_o;
  wire _al_u5705_o;
  wire _al_u5706_o;
  wire _al_u5707_o;
  wire _al_u5708_o;
  wire _al_u5709_o;
  wire _al_u5710_o;
  wire _al_u5711_o;
  wire _al_u5712_o;
  wire _al_u5713_o;
  wire _al_u5714_o;
  wire _al_u5715_o;
  wire _al_u5716_o;
  wire _al_u5717_o;
  wire _al_u5718_o;
  wire _al_u5719_o;
  wire _al_u571_o;
  wire _al_u5720_o;
  wire _al_u5721_o;
  wire _al_u5722_o;
  wire _al_u5723_o;
  wire _al_u5724_o;
  wire _al_u5725_o;
  wire _al_u5726_o;
  wire _al_u5727_o;
  wire _al_u5728_o;
  wire _al_u5729_o;
  wire _al_u572_o;
  wire _al_u5730_o;
  wire _al_u5731_o;
  wire _al_u5732_o;
  wire _al_u5733_o;
  wire _al_u5734_o;
  wire _al_u5735_o;
  wire _al_u5736_o;
  wire _al_u5737_o;
  wire _al_u5738_o;
  wire _al_u5739_o;
  wire _al_u573_o;
  wire _al_u5740_o;
  wire _al_u5741_o;
  wire _al_u5742_o;
  wire _al_u5743_o;
  wire _al_u5744_o;
  wire _al_u5745_o;
  wire _al_u5746_o;
  wire _al_u5747_o;
  wire _al_u5748_o;
  wire _al_u5749_o;
  wire _al_u574_o;
  wire _al_u5750_o;
  wire _al_u5751_o;
  wire _al_u5752_o;
  wire _al_u5753_o;
  wire _al_u5754_o;
  wire _al_u5755_o;
  wire _al_u5756_o;
  wire _al_u5757_o;
  wire _al_u5758_o;
  wire _al_u5759_o;
  wire _al_u575_o;
  wire _al_u5760_o;
  wire _al_u5761_o;
  wire _al_u5762_o;
  wire _al_u5763_o;
  wire _al_u5764_o;
  wire _al_u5765_o;
  wire _al_u5766_o;
  wire _al_u5767_o;
  wire _al_u5768_o;
  wire _al_u5769_o;
  wire _al_u576_o;
  wire _al_u5770_o;
  wire _al_u5771_o;
  wire _al_u5772_o;
  wire _al_u5773_o;
  wire _al_u5774_o;
  wire _al_u5775_o;
  wire _al_u5776_o;
  wire _al_u5777_o;
  wire _al_u5778_o;
  wire _al_u5779_o;
  wire _al_u5780_o;
  wire _al_u5782_o;
  wire _al_u5783_o;
  wire _al_u5784_o;
  wire _al_u5785_o;
  wire _al_u5786_o;
  wire _al_u5787_o;
  wire _al_u5788_o;
  wire _al_u5789_o;
  wire _al_u5790_o;
  wire _al_u5791_o;
  wire _al_u5792_o;
  wire _al_u5793_o;
  wire _al_u5794_o;
  wire _al_u5795_o;
  wire _al_u5796_o;
  wire _al_u5797_o;
  wire _al_u5798_o;
  wire _al_u5799_o;
  wire _al_u5800_o;
  wire _al_u5801_o;
  wire _al_u5802_o;
  wire _al_u5803_o;
  wire _al_u5804_o;
  wire _al_u5805_o;
  wire _al_u5806_o;
  wire _al_u5807_o;
  wire _al_u5808_o;
  wire _al_u5809_o;
  wire _al_u580_o;
  wire _al_u5810_o;
  wire _al_u5812_o;
  wire _al_u5813_o;
  wire _al_u5814_o;
  wire _al_u5816_o;
  wire _al_u5818_o;
  wire _al_u581_o;
  wire _al_u5820_o;
  wire _al_u5822_o;
  wire _al_u5824_o;
  wire _al_u5826_o;
  wire _al_u5828_o;
  wire _al_u582_o;
  wire _al_u5830_o;
  wire _al_u5832_o;
  wire _al_u5834_o;
  wire _al_u5836_o;
  wire _al_u5843_o;
  wire _al_u5845_o;
  wire _al_u5848_o;
  wire _al_u584_o;
  wire _al_u5850_o;
  wire _al_u5851_o;
  wire _al_u5853_o;
  wire _al_u5854_o;
  wire _al_u5856_o;
  wire _al_u5857_o;
  wire _al_u5858_o;
  wire _al_u5859_o;
  wire _al_u585_o;
  wire _al_u5860_o;
  wire _al_u5861_o;
  wire _al_u5862_o;
  wire _al_u5864_o;
  wire _al_u5865_o;
  wire _al_u5866_o;
  wire _al_u5868_o;
  wire _al_u5869_o;
  wire _al_u5870_o;
  wire _al_u5871_o;
  wire _al_u5872_o;
  wire _al_u5873_o;
  wire _al_u5874_o;
  wire _al_u5875_o;
  wire _al_u5878_o;
  wire _al_u5879_o;
  wire _al_u587_o;
  wire _al_u5880_o;
  wire _al_u5883_o;
  wire _al_u5884_o;
  wire _al_u5885_o;
  wire _al_u5886_o;
  wire _al_u5887_o;
  wire _al_u5888_o;
  wire _al_u5889_o;
  wire _al_u588_o;
  wire _al_u5890_o;
  wire _al_u5891_o;
  wire _al_u5892_o;
  wire _al_u5893_o;
  wire _al_u5894_o;
  wire _al_u5896_o;
  wire _al_u5897_o;
  wire _al_u5899_o;
  wire _al_u5900_o;
  wire _al_u5903_o;
  wire _al_u5904_o;
  wire _al_u5905_o;
  wire _al_u5906_o;
  wire _al_u5908_o;
  wire _al_u5909_o;
  wire _al_u5910_o;
  wire _al_u5911_o;
  wire _al_u5912_o;
  wire _al_u5913_o;
  wire _al_u5915_o;
  wire _al_u5916_o;
  wire _al_u5917_o;
  wire _al_u5918_o;
  wire _al_u5919_o;
  wire _al_u591_o;
  wire _al_u5920_o;
  wire _al_u5921_o;
  wire _al_u5922_o;
  wire _al_u5924_o;
  wire _al_u5925_o;
  wire _al_u5926_o;
  wire _al_u5927_o;
  wire _al_u5929_o;
  wire _al_u5930_o;
  wire _al_u5931_o;
  wire _al_u5932_o;
  wire _al_u5933_o;
  wire _al_u5934_o;
  wire _al_u5935_o;
  wire _al_u5936_o;
  wire _al_u5937_o;
  wire _al_u5938_o;
  wire _al_u593_o;
  wire _al_u5940_o;
  wire _al_u5941_o;
  wire _al_u5942_o;
  wire _al_u5943_o;
  wire _al_u5945_o;
  wire _al_u5946_o;
  wire _al_u5947_o;
  wire _al_u5948_o;
  wire _al_u5950_o;
  wire _al_u5951_o;
  wire _al_u5952_o;
  wire _al_u5953_o;
  wire _al_u5954_o;
  wire _al_u5955_o;
  wire _al_u5956_o;
  wire _al_u5957_o;
  wire _al_u5958_o;
  wire _al_u5959_o;
  wire _al_u5960_o;
  wire _al_u5961_o;
  wire _al_u5963_o;
  wire _al_u5964_o;
  wire _al_u5966_o;
  wire _al_u5968_o;
  wire _al_u5969_o;
  wire _al_u5970_o;
  wire _al_u5971_o;
  wire _al_u5972_o;
  wire _al_u5973_o;
  wire _al_u5974_o;
  wire _al_u5977_o;
  wire _al_u5979_o;
  wire _al_u597_o;
  wire _al_u5980_o;
  wire _al_u5983_o;
  wire _al_u5984_o;
  wire _al_u5985_o;
  wire _al_u5987_o;
  wire _al_u5988_o;
  wire _al_u5990_o;
  wire _al_u5991_o;
  wire _al_u5993_o;
  wire _al_u5995_o;
  wire _al_u5998_o;
  wire _al_u6000_o;
  wire _al_u6002_o;
  wire _al_u6003_o;
  wire _al_u6004_o;
  wire _al_u6005_o;
  wire _al_u6006_o;
  wire _al_u6007_o;
  wire _al_u6008_o;
  wire _al_u6009_o;
  wire _al_u6010_o;
  wire _al_u6011_o;
  wire _al_u6013_o;
  wire _al_u6014_o;
  wire _al_u6015_o;
  wire _al_u6016_o;
  wire _al_u6017_o;
  wire _al_u6018_o;
  wire _al_u6021_o;
  wire _al_u6023_o;
  wire _al_u6024_o;
  wire _al_u6025_o;
  wire _al_u6026_o;
  wire _al_u6027_o;
  wire _al_u6028_o;
  wire _al_u6029_o;
  wire _al_u6030_o;
  wire _al_u6032_o;
  wire _al_u6033_o;
  wire _al_u6034_o;
  wire _al_u6035_o;
  wire _al_u6036_o;
  wire _al_u6037_o;
  wire _al_u6039_o;
  wire _al_u6040_o;
  wire _al_u6041_o;
  wire _al_u6042_o;
  wire _al_u6043_o;
  wire _al_u6044_o;
  wire _al_u6045_o;
  wire _al_u6046_o;
  wire _al_u6047_o;
  wire _al_u6049_o;
  wire _al_u604_o;
  wire _al_u6050_o;
  wire _al_u6052_o;
  wire _al_u6053_o;
  wire _al_u6054_o;
  wire _al_u6055_o;
  wire _al_u6056_o;
  wire _al_u6057_o;
  wire _al_u6059_o;
  wire _al_u6060_o;
  wire _al_u6061_o;
  wire _al_u6062_o;
  wire _al_u6063_o;
  wire _al_u6064_o;
  wire _al_u6065_o;
  wire _al_u6066_o;
  wire _al_u6067_o;
  wire _al_u6068_o;
  wire _al_u6069_o;
  wire _al_u606_o;
  wire _al_u6070_o;
  wire _al_u6071_o;
  wire _al_u6073_o;
  wire _al_u6074_o;
  wire _al_u6075_o;
  wire _al_u6076_o;
  wire _al_u6077_o;
  wire _al_u6078_o;
  wire _al_u6079_o;
  wire _al_u607_o;
  wire _al_u6080_o;
  wire _al_u6081_o;
  wire _al_u6082_o;
  wire _al_u6084_o;
  wire _al_u6085_o;
  wire _al_u6086_o;
  wire _al_u6087_o;
  wire _al_u6088_o;
  wire _al_u6089_o;
  wire _al_u6091_o;
  wire _al_u6092_o;
  wire _al_u6094_o;
  wire _al_u6095_o;
  wire _al_u6096_o;
  wire _al_u6099_o;
  wire _al_u609_o;
  wire _al_u6100_o;
  wire _al_u6101_o;
  wire _al_u6102_o;
  wire _al_u6103_o;
  wire _al_u6104_o;
  wire _al_u6105_o;
  wire _al_u6106_o;
  wire _al_u6108_o;
  wire _al_u6109_o;
  wire _al_u6112_o;
  wire _al_u6113_o;
  wire _al_u6115_o;
  wire _al_u6116_o;
  wire _al_u6118_o;
  wire _al_u6120_o;
  wire _al_u6121_o;
  wire _al_u6122_o;
  wire _al_u6123_o;
  wire _al_u6124_o;
  wire _al_u6125_o;
  wire _al_u6127_o;
  wire _al_u6128_o;
  wire _al_u6129_o;
  wire _al_u6130_o;
  wire _al_u6133_o;
  wire _al_u6134_o;
  wire _al_u6135_o;
  wire _al_u6137_o;
  wire _al_u6138_o;
  wire _al_u6139_o;
  wire _al_u6141_o;
  wire _al_u6142_o;
  wire _al_u6144_o;
  wire _al_u6145_o;
  wire _al_u6147_o;
  wire _al_u6149_o;
  wire _al_u6150_o;
  wire _al_u6151_o;
  wire _al_u6153_o;
  wire _al_u6154_o;
  wire _al_u6155_o;
  wire _al_u6157_o;
  wire _al_u6158_o;
  wire _al_u6159_o;
  wire _al_u6160_o;
  wire _al_u6161_o;
  wire _al_u6163_o;
  wire _al_u6164_o;
  wire _al_u6166_o;
  wire _al_u6167_o;
  wire _al_u6168_o;
  wire _al_u6169_o;
  wire _al_u6170_o;
  wire _al_u6171_o;
  wire _al_u6172_o;
  wire _al_u6173_o;
  wire _al_u6174_o;
  wire _al_u6175_o;
  wire _al_u6176_o;
  wire _al_u6177_o;
  wire _al_u6180_o;
  wire _al_u6181_o;
  wire _al_u6182_o;
  wire _al_u6183_o;
  wire _al_u6184_o;
  wire _al_u6185_o;
  wire _al_u6186_o;
  wire _al_u6187_o;
  wire _al_u6188_o;
  wire _al_u6189_o;
  wire _al_u6190_o;
  wire _al_u6191_o;
  wire _al_u6192_o;
  wire _al_u6193_o;
  wire _al_u6194_o;
  wire _al_u6196_o;
  wire _al_u6197_o;
  wire _al_u6198_o;
  wire _al_u6200_o;
  wire _al_u6201_o;
  wire _al_u6202_o;
  wire _al_u6203_o;
  wire _al_u6205_o;
  wire _al_u6206_o;
  wire _al_u6207_o;
  wire _al_u6208_o;
  wire _al_u6210_o;
  wire _al_u6211_o;
  wire _al_u6214_o;
  wire _al_u6216_o;
  wire _al_u6217_o;
  wire _al_u6218_o;
  wire _al_u6219_o;
  wire _al_u6220_o;
  wire _al_u6222_o;
  wire _al_u6225_o;
  wire _al_u6226_o;
  wire _al_u6227_o;
  wire _al_u6228_o;
  wire _al_u6229_o;
  wire _al_u6230_o;
  wire _al_u6231_o;
  wire _al_u6232_o;
  wire _al_u6233_o;
  wire _al_u6234_o;
  wire _al_u6235_o;
  wire _al_u6236_o;
  wire _al_u6237_o;
  wire _al_u6238_o;
  wire _al_u6240_o;
  wire _al_u6241_o;
  wire _al_u6242_o;
  wire _al_u6243_o;
  wire _al_u6244_o;
  wire _al_u6246_o;
  wire _al_u6248_o;
  wire _al_u6249_o;
  wire _al_u6251_o;
  wire _al_u6252_o;
  wire _al_u6253_o;
  wire _al_u6254_o;
  wire _al_u6255_o;
  wire _al_u6256_o;
  wire _al_u6257_o;
  wire _al_u6258_o;
  wire _al_u6259_o;
  wire _al_u6260_o;
  wire _al_u6261_o;
  wire _al_u6262_o;
  wire _al_u6263_o;
  wire _al_u6264_o;
  wire _al_u6265_o;
  wire _al_u6266_o;
  wire _al_u6267_o;
  wire _al_u6268_o;
  wire _al_u6269_o;
  wire _al_u6271_o;
  wire _al_u6273_o;
  wire _al_u6274_o;
  wire _al_u6275_o;
  wire _al_u6276_o;
  wire _al_u6277_o;
  wire _al_u6278_o;
  wire _al_u6279_o;
  wire _al_u6280_o;
  wire _al_u6281_o;
  wire _al_u6284_o;
  wire _al_u6285_o;
  wire _al_u6286_o;
  wire _al_u6287_o;
  wire _al_u6288_o;
  wire _al_u6289_o;
  wire _al_u6290_o;
  wire _al_u6291_o;
  wire _al_u6292_o;
  wire _al_u6293_o;
  wire _al_u6294_o;
  wire _al_u6295_o;
  wire _al_u6296_o;
  wire _al_u6298_o;
  wire _al_u6300_o;
  wire _al_u6302_o;
  wire _al_u6304_o;
  wire _al_u6306_o;
  wire _al_u6307_o;
  wire _al_u6308_o;
  wire _al_u6310_o;
  wire _al_u6311_o;
  wire _al_u6312_o;
  wire _al_u6313_o;
  wire _al_u6314_o;
  wire _al_u6315_o;
  wire _al_u6316_o;
  wire _al_u6317_o;
  wire _al_u6318_o;
  wire _al_u6319_o;
  wire _al_u6320_o;
  wire _al_u6321_o;
  wire _al_u6322_o;
  wire _al_u6323_o;
  wire _al_u6324_o;
  wire _al_u6325_o;
  wire _al_u6326_o;
  wire _al_u6327_o;
  wire _al_u6328_o;
  wire _al_u6329_o;
  wire _al_u6331_o;
  wire _al_u6332_o;
  wire _al_u6333_o;
  wire _al_u6335_o;
  wire _al_u6336_o;
  wire _al_u6337_o;
  wire _al_u6338_o;
  wire _al_u6339_o;
  wire _al_u6341_o;
  wire _al_u6342_o;
  wire _al_u6343_o;
  wire _al_u6344_o;
  wire _al_u6345_o;
  wire _al_u6347_o;
  wire _al_u6348_o;
  wire _al_u6349_o;
  wire _al_u6350_o;
  wire _al_u6351_o;
  wire _al_u6352_o;
  wire _al_u6353_o;
  wire _al_u6354_o;
  wire _al_u6355_o;
  wire _al_u6356_o;
  wire _al_u6357_o;
  wire _al_u6358_o;
  wire _al_u6360_o;
  wire _al_u6361_o;
  wire _al_u6362_o;
  wire _al_u6363_o;
  wire _al_u6364_o;
  wire _al_u6365_o;
  wire _al_u6367_o;
  wire _al_u6368_o;
  wire _al_u6369_o;
  wire _al_u6370_o;
  wire _al_u6371_o;
  wire _al_u6372_o;
  wire _al_u6373_o;
  wire _al_u637_o;
  wire _al_u6380_o;
  wire _al_u6381_o;
  wire _al_u6382_o;
  wire _al_u6383_o;
  wire _al_u6384_o;
  wire _al_u6385_o;
  wire _al_u6388_o;
  wire _al_u6389_o;
  wire _al_u6390_o;
  wire _al_u6392_o;
  wire _al_u6393_o;
  wire _al_u6394_o;
  wire _al_u6395_o;
  wire _al_u6396_o;
  wire _al_u6397_o;
  wire _al_u6398_o;
  wire _al_u6399_o;
  wire _al_u6400_o;
  wire _al_u6401_o;
  wire _al_u6402_o;
  wire _al_u6403_o;
  wire _al_u6404_o;
  wire _al_u6405_o;
  wire _al_u6406_o;
  wire _al_u6407_o;
  wire _al_u6408_o;
  wire _al_u6409_o;
  wire _al_u6410_o;
  wire _al_u6411_o;
  wire _al_u6412_o;
  wire _al_u6413_o;
  wire _al_u6416_o;
  wire _al_u6417_o;
  wire _al_u6418_o;
  wire _al_u6419_o;
  wire _al_u6420_o;
  wire _al_u6421_o;
  wire _al_u6422_o;
  wire _al_u6423_o;
  wire _al_u6431_o;
  wire _al_u6432_o;
  wire _al_u6433_o;
  wire _al_u6434_o;
  wire _al_u6435_o;
  wire _al_u6436_o;
  wire _al_u6437_o;
  wire _al_u6438_o;
  wire _al_u6439_o;
  wire _al_u6440_o;
  wire _al_u6441_o;
  wire _al_u6442_o;
  wire _al_u6443_o;
  wire _al_u6444_o;
  wire _al_u6446_o;
  wire _al_u6447_o;
  wire _al_u6448_o;
  wire _al_u6449_o;
  wire _al_u6450_o;
  wire _al_u6451_o;
  wire _al_u6452_o;
  wire _al_u6453_o;
  wire _al_u6454_o;
  wire _al_u6455_o;
  wire _al_u6457_o;
  wire _al_u6458_o;
  wire _al_u6459_o;
  wire _al_u6460_o;
  wire _al_u6461_o;
  wire _al_u6463_o;
  wire _al_u6464_o;
  wire _al_u6467_o;
  wire _al_u6468_o;
  wire _al_u6469_o;
  wire _al_u6471_o;
  wire _al_u6472_o;
  wire _al_u6473_o;
  wire _al_u6475_o;
  wire _al_u6476_o;
  wire _al_u6477_o;
  wire _al_u6478_o;
  wire _al_u6479_o;
  wire _al_u6480_o;
  wire _al_u6481_o;
  wire _al_u6482_o;
  wire _al_u6483_o;
  wire _al_u6484_o;
  wire _al_u6491_o;
  wire _al_u6492_o;
  wire _al_u6493_o;
  wire _al_u6494_o;
  wire _al_u6495_o;
  wire _al_u6497_o;
  wire _al_u6498_o;
  wire _al_u6499_o;
  wire _al_u6500_o;
  wire _al_u6501_o;
  wire _al_u6502_o;
  wire _al_u6503_o;
  wire _al_u6504_o;
  wire _al_u6505_o;
  wire _al_u6507_o;
  wire _al_u6508_o;
  wire _al_u6509_o;
  wire _al_u650_o;
  wire _al_u6510_o;
  wire _al_u6511_o;
  wire _al_u6512_o;
  wire _al_u6513_o;
  wire _al_u6515_o;
  wire _al_u6518_o;
  wire _al_u6519_o;
  wire _al_u6520_o;
  wire _al_u6521_o;
  wire _al_u6522_o;
  wire _al_u6524_o;
  wire _al_u6525_o;
  wire _al_u6526_o;
  wire _al_u6527_o;
  wire _al_u6528_o;
  wire _al_u6529_o;
  wire _al_u6530_o;
  wire _al_u6531_o;
  wire _al_u6532_o;
  wire _al_u6533_o;
  wire _al_u6534_o;
  wire _al_u6535_o;
  wire _al_u6538_o;
  wire _al_u6540_o;
  wire _al_u6541_o;
  wire _al_u6542_o;
  wire _al_u6543_o;
  wire _al_u6544_o;
  wire _al_u6545_o;
  wire _al_u6546_o;
  wire _al_u6547_o;
  wire _al_u6548_o;
  wire _al_u6549_o;
  wire _al_u6550_o;
  wire _al_u6551_o;
  wire _al_u6552_o;
  wire _al_u6553_o;
  wire _al_u6554_o;
  wire _al_u6555_o;
  wire _al_u6556_o;
  wire _al_u6557_o;
  wire _al_u6558_o;
  wire _al_u6560_o;
  wire _al_u6562_o;
  wire _al_u6563_o;
  wire _al_u6564_o;
  wire _al_u6565_o;
  wire _al_u6566_o;
  wire _al_u6567_o;
  wire _al_u6568_o;
  wire _al_u6569_o;
  wire _al_u6570_o;
  wire _al_u6571_o;
  wire _al_u6572_o;
  wire _al_u6573_o;
  wire _al_u6574_o;
  wire _al_u6575_o;
  wire _al_u6576_o;
  wire _al_u6577_o;
  wire _al_u6578_o;
  wire _al_u6579_o;
  wire _al_u6580_o;
  wire _al_u6581_o;
  wire _al_u6582_o;
  wire _al_u6583_o;
  wire _al_u6584_o;
  wire _al_u6586_o;
  wire _al_u6587_o;
  wire _al_u6588_o;
  wire _al_u6589_o;
  wire _al_u6590_o;
  wire _al_u6591_o;
  wire _al_u6592_o;
  wire _al_u6593_o;
  wire _al_u6596_o;
  wire _al_u6599_o;
  wire _al_u6600_o;
  wire _al_u6601_o;
  wire _al_u6602_o;
  wire _al_u6603_o;
  wire _al_u6604_o;
  wire _al_u6605_o;
  wire _al_u6610_o;
  wire _al_u6611_o;
  wire _al_u6612_o;
  wire _al_u6614_o;
  wire _al_u6615_o;
  wire _al_u6616_o;
  wire _al_u6617_o;
  wire _al_u6619_o;
  wire _al_u6620_o;
  wire _al_u6621_o;
  wire _al_u6624_o;
  wire _al_u6625_o;
  wire _al_u6626_o;
  wire _al_u6627_o;
  wire _al_u6628_o;
  wire _al_u6629_o;
  wire _al_u6631_o;
  wire _al_u6632_o;
  wire _al_u6633_o;
  wire _al_u6634_o;
  wire _al_u6635_o;
  wire _al_u6636_o;
  wire _al_u6637_o;
  wire _al_u6638_o;
  wire _al_u6639_o;
  wire _al_u6640_o;
  wire _al_u6641_o;
  wire _al_u6643_o;
  wire _al_u6645_o;
  wire _al_u6646_o;
  wire _al_u6647_o;
  wire _al_u6648_o;
  wire _al_u6649_o;
  wire _al_u6650_o;
  wire _al_u6651_o;
  wire _al_u6652_o;
  wire _al_u6653_o;
  wire _al_u6654_o;
  wire _al_u6655_o;
  wire _al_u6656_o;
  wire _al_u6658_o;
  wire _al_u6659_o;
  wire _al_u6660_o;
  wire _al_u6661_o;
  wire _al_u6662_o;
  wire _al_u6663_o;
  wire _al_u6664_o;
  wire _al_u6665_o;
  wire _al_u6666_o;
  wire _al_u6667_o;
  wire _al_u6668_o;
  wire _al_u6669_o;
  wire _al_u6670_o;
  wire _al_u6672_o;
  wire _al_u6673_o;
  wire _al_u6674_o;
  wire _al_u6675_o;
  wire _al_u6676_o;
  wire _al_u6677_o;
  wire _al_u6679_o;
  wire _al_u6680_o;
  wire _al_u6681_o;
  wire _al_u6682_o;
  wire _al_u6683_o;
  wire _al_u6684_o;
  wire _al_u6686_o;
  wire _al_u6687_o;
  wire _al_u6688_o;
  wire _al_u6689_o;
  wire _al_u6690_o;
  wire _al_u6691_o;
  wire _al_u6692_o;
  wire _al_u6693_o;
  wire _al_u6694_o;
  wire _al_u6695_o;
  wire _al_u6696_o;
  wire _al_u6697_o;
  wire _al_u6698_o;
  wire _al_u6699_o;
  wire _al_u6700_o;
  wire _al_u6701_o;
  wire _al_u6702_o;
  wire _al_u6703_o;
  wire _al_u6706_o;
  wire _al_u6708_o;
  wire _al_u6709_o;
  wire _al_u6710_o;
  wire _al_u6711_o;
  wire _al_u6712_o;
  wire _al_u6713_o;
  wire _al_u6714_o;
  wire _al_u6715_o;
  wire _al_u6716_o;
  wire _al_u6717_o;
  wire _al_u6718_o;
  wire _al_u6719_o;
  wire _al_u6720_o;
  wire _al_u6721_o;
  wire _al_u6722_o;
  wire _al_u6723_o;
  wire _al_u6724_o;
  wire _al_u6725_o;
  wire _al_u6727_o;
  wire _al_u6728_o;
  wire _al_u6729_o;
  wire _al_u6730_o;
  wire _al_u6731_o;
  wire _al_u6732_o;
  wire _al_u6733_o;
  wire _al_u6734_o;
  wire _al_u6735_o;
  wire _al_u6737_o;
  wire _al_u6738_o;
  wire _al_u6740_o;
  wire _al_u6741_o;
  wire _al_u6742_o;
  wire _al_u6743_o;
  wire _al_u6744_o;
  wire _al_u6745_o;
  wire _al_u6746_o;
  wire _al_u6749_o;
  wire _al_u6751_o;
  wire _al_u6752_o;
  wire _al_u6753_o;
  wire _al_u6754_o;
  wire _al_u6755_o;
  wire _al_u6756_o;
  wire _al_u6757_o;
  wire _al_u6758_o;
  wire _al_u6759_o;
  wire _al_u6760_o;
  wire _al_u6761_o;
  wire _al_u6762_o;
  wire _al_u6765_o;
  wire _al_u6767_o;
  wire _al_u6769_o;
  wire _al_u6771_o;
  wire _al_u6773_o;
  wire _al_u6775_o;
  wire _al_u6776_o;
  wire _al_u6778_o;
  wire _al_u677_o;
  wire _al_u6780_o;
  wire _al_u6782_o;
  wire _al_u6784_o;
  wire _al_u6786_o;
  wire _al_u6788_o;
  wire _al_u678_o;
  wire _al_u6790_o;
  wire _al_u6792_o;
  wire _al_u6794_o;
  wire _al_u6795_o;
  wire _al_u6796_o;
  wire _al_u6797_o;
  wire _al_u6798_o;
  wire _al_u6799_o;
  wire _al_u679_o;
  wire _al_u6800_o;
  wire _al_u6801_o;
  wire _al_u6802_o;
  wire _al_u6803_o;
  wire _al_u6805_o;
  wire _al_u6806_o;
  wire _al_u6807_o;
  wire _al_u6808_o;
  wire _al_u6809_o;
  wire _al_u680_o;
  wire _al_u6810_o;
  wire _al_u6811_o;
  wire _al_u6812_o;
  wire _al_u6814_o;
  wire _al_u6817_o;
  wire _al_u6819_o;
  wire _al_u681_o;
  wire _al_u6820_o;
  wire _al_u6821_o;
  wire _al_u6822_o;
  wire _al_u6823_o;
  wire _al_u6824_o;
  wire _al_u6825_o;
  wire _al_u6826_o;
  wire _al_u6827_o;
  wire _al_u6828_o;
  wire _al_u6829_o;
  wire _al_u682_o;
  wire _al_u6830_o;
  wire _al_u6832_o;
  wire _al_u6833_o;
  wire _al_u6836_o;
  wire _al_u6838_o;
  wire _al_u6841_o;
  wire _al_u6842_o;
  wire _al_u6844_o;
  wire _al_u6846_o;
  wire _al_u6848_o;
  wire _al_u6850_o;
  wire _al_u6852_o;
  wire _al_u6853_o;
  wire _al_u6855_o;
  wire _al_u6856_o;
  wire _al_u6857_o;
  wire _al_u6858_o;
  wire _al_u6859_o;
  wire _al_u685_o;
  wire _al_u6861_o;
  wire _al_u6866_o;
  wire _al_u6867_o;
  wire _al_u6868_o;
  wire _al_u6869_o;
  wire _al_u6870_o;
  wire _al_u6871_o;
  wire _al_u6872_o;
  wire _al_u6874_o;
  wire _al_u6875_o;
  wire _al_u6876_o;
  wire _al_u6878_o;
  wire _al_u6879_o;
  wire _al_u6881_o;
  wire _al_u6882_o;
  wire _al_u6884_o;
  wire _al_u6885_o;
  wire _al_u6887_o;
  wire _al_u6888_o;
  wire _al_u6890_o;
  wire _al_u6891_o;
  wire _al_u6892_o;
  wire _al_u6894_o;
  wire _al_u6897_o;
  wire _al_u6898_o;
  wire _al_u6900_o;
  wire _al_u6901_o;
  wire _al_u6903_o;
  wire _al_u6904_o;
  wire _al_u6907_o;
  wire _al_u6908_o;
  wire _al_u6910_o;
  wire _al_u6913_o;
  wire _al_u6914_o;
  wire _al_u6915_o;
  wire _al_u6917_o;
  wire _al_u6918_o;
  wire _al_u6920_o;
  wire _al_u6921_o;
  wire _al_u6923_o;
  wire _al_u6924_o;
  wire _al_u6925_o;
  wire _al_u6926_o;
  wire _al_u6929_o;
  wire _al_u692_o;
  wire _al_u6930_o;
  wire _al_u6931_o;
  wire _al_u6932_o;
  wire _al_u6934_o;
  wire _al_u6935_o;
  wire _al_u6937_o;
  wire _al_u6938_o;
  wire _al_u6941_o;
  wire _al_u6942_o;
  wire _al_u6945_o;
  wire _al_u6946_o;
  wire _al_u6947_o;
  wire _al_u6948_o;
  wire _al_u6949_o;
  wire _al_u6950_o;
  wire _al_u6951_o;
  wire _al_u6952_o;
  wire _al_u6953_o;
  wire _al_u6954_o;
  wire _al_u6956_o;
  wire _al_u6957_o;
  wire _al_u6958_o;
  wire _al_u695_o;
  wire _al_u6960_o;
  wire _al_u6961_o;
  wire _al_u6962_o;
  wire _al_u6964_o;
  wire _al_u6965_o;
  wire _al_u6966_o;
  wire _al_u6967_o;
  wire _al_u6968_o;
  wire _al_u6969_o;
  wire _al_u696_o;
  wire _al_u6970_o;
  wire _al_u6972_o;
  wire _al_u6975_o;
  wire _al_u6977_o;
  wire _al_u6978_o;
  wire _al_u6979_o;
  wire _al_u697_o;
  wire _al_u6980_o;
  wire _al_u6981_o;
  wire _al_u6983_o;
  wire _al_u6984_o;
  wire _al_u6985_o;
  wire _al_u6987_o;
  wire _al_u6988_o;
  wire _al_u6989_o;
  wire _al_u698_o;
  wire _al_u6992_o;
  wire _al_u6993_o;
  wire _al_u6994_o;
  wire _al_u6996_o;
  wire _al_u6997_o;
  wire _al_u6998_o;
  wire _al_u7000_o;
  wire _al_u7001_o;
  wire _al_u7002_o;
  wire _al_u7005_o;
  wire _al_u7006_o;
  wire _al_u7008_o;
  wire _al_u7009_o;
  wire _al_u700_o;
  wire _al_u7010_o;
  wire _al_u7012_o;
  wire _al_u7013_o;
  wire _al_u7014_o;
  wire _al_u7015_o;
  wire _al_u7016_o;
  wire _al_u7018_o;
  wire _al_u7020_o;
  wire _al_u7021_o;
  wire _al_u7022_o;
  wire _al_u7023_o;
  wire _al_u7024_o;
  wire _al_u7025_o;
  wire _al_u7027_o;
  wire _al_u7028_o;
  wire _al_u702_o;
  wire _al_u7030_o;
  wire _al_u7031_o;
  wire _al_u7032_o;
  wire _al_u7034_o;
  wire _al_u7035_o;
  wire _al_u7036_o;
  wire _al_u7038_o;
  wire _al_u7039_o;
  wire _al_u7040_o;
  wire _al_u7041_o;
  wire _al_u7044_o;
  wire _al_u7045_o;
  wire _al_u7047_o;
  wire _al_u7048_o;
  wire _al_u7049_o;
  wire _al_u7051_o;
  wire _al_u7052_o;
  wire _al_u7053_o;
  wire _al_u7056_o;
  wire _al_u7057_o;
  wire _al_u7059_o;
  wire _al_u705_o;
  wire _al_u7060_o;
  wire _al_u7062_o;
  wire _al_u7064_o;
  wire _al_u7065_o;
  wire _al_u7068_o;
  wire _al_u7069_o;
  wire _al_u7071_o;
  wire _al_u7072_o;
  wire _al_u7074_o;
  wire _al_u7075_o;
  wire _al_u7077_o;
  wire _al_u7078_o;
  wire _al_u7080_o;
  wire _al_u7081_o;
  wire _al_u7083_o;
  wire _al_u7084_o;
  wire _al_u7085_o;
  wire _al_u7087_o;
  wire _al_u7088_o;
  wire _al_u7090_o;
  wire _al_u7092_o;
  wire _al_u7093_o;
  wire _al_u7094_o;
  wire _al_u7096_o;
  wire _al_u7097_o;
  wire _al_u7099_o;
  wire _al_u7100_o;
  wire _al_u7101_o;
  wire _al_u7103_o;
  wire _al_u7104_o;
  wire _al_u7105_o;
  wire _al_u7108_o;
  wire _al_u7109_o;
  wire _al_u7112_o;
  wire _al_u7113_o;
  wire _al_u7116_o;
  wire _al_u7117_o;
  wire _al_u7119_o;
  wire _al_u711_o;
  wire _al_u7120_o;
  wire _al_u7121_o;
  wire _al_u7122_o;
  wire _al_u7124_o;
  wire _al_u7125_o;
  wire _al_u7126_o;
  wire _al_u7128_o;
  wire _al_u7130_o;
  wire _al_u7131_o;
  wire _al_u7133_o;
  wire _al_u7135_o;
  wire _al_u7137_o;
  wire _al_u7139_o;
  wire _al_u7141_o;
  wire _al_u7144_o;
  wire _al_u7146_o;
  wire _al_u7148_o;
  wire _al_u714_o;
  wire _al_u7151_o;
  wire _al_u7154_o;
  wire _al_u7157_o;
  wire _al_u7160_o;
  wire _al_u7163_o;
  wire _al_u7166_o;
  wire _al_u7169_o;
  wire _al_u7172_o;
  wire _al_u7175_o;
  wire _al_u7178_o;
  wire _al_u717_o;
  wire _al_u7181_o;
  wire _al_u7184_o;
  wire _al_u7187_o;
  wire _al_u718_o;
  wire _al_u7190_o;
  wire _al_u7193_o;
  wire _al_u7195_o;
  wire _al_u7198_o;
  wire _al_u719_o;
  wire _al_u7201_o;
  wire _al_u7204_o;
  wire _al_u7206_o;
  wire _al_u7207_o;
  wire _al_u7208_o;
  wire _al_u720_o;
  wire _al_u7211_o;
  wire _al_u7214_o;
  wire _al_u7217_o;
  wire _al_u7220_o;
  wire _al_u7222_o;
  wire _al_u7223_o;
  wire _al_u7224_o;
  wire _al_u7225_o;
  wire _al_u723_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u729_o;
  wire _al_u731_o;
  wire _al_u732_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u744_o;
  wire _al_u747_o;
  wire _al_u749_o;
  wire _al_u750_o;
  wire _al_u753_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u759_o;
  wire _al_u760_o;
  wire _al_u761_o;
  wire _al_u762_o;
  wire _al_u765_o;
  wire _al_u766_o;
  wire _al_u767_o;
  wire _al_u768_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u774_o;
  wire _al_u777_o;
  wire _al_u778_o;
  wire _al_u779_o;
  wire _al_u780_o;
  wire _al_u783_o;
  wire _al_u786_o;
  wire _al_u789_o;
  wire _al_u790_o;
  wire _al_u792_o;
  wire _al_u795_o;
  wire _al_u796_o;
  wire _al_u797_o;
  wire _al_u798_o;
  wire _al_u801_o;
  wire _al_u802_o;
  wire _al_u804_o;
  wire _al_u807_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u815_o;
  wire _al_u816_o;
  wire _al_u819_o;
  wire _al_u821_o;
  wire _al_u822_o;
  wire _al_u823_o;
  wire _al_u825_o;
  wire _al_u828_o;
  wire _al_u831_o;
  wire _al_u832_o;
  wire _al_u833_o;
  wire _al_u837_o;
  wire _al_u839_o;
  wire _al_u840_o;
  wire _al_u843_o;
  wire _al_u844_o;
  wire _al_u846_o;
  wire _al_u849_o;
  wire _al_u850_o;
  wire _al_u851_o;
  wire _al_u852_o;
  wire _al_u855_o;
  wire _al_u858_o;
  wire _al_u861_o;
  wire _al_u862_o;
  wire _al_u864_o;
  wire _al_u867_o;
  wire _al_u868_o;
  wire _al_u869_o;
  wire _al_u870_o;
  wire _al_u873_o;
  wire _al_u874_o;
  wire _al_u875_o;
  wire _al_u876_o;
  wire _al_u879_o;
  wire _al_u880_o;
  wire _al_u882_o;
  wire _al_u885_o;
  wire _al_u886_o;
  wire _al_u887_o;
  wire _al_u888_o;
  wire _al_u891_o;
  wire _al_u892_o;
  wire _al_u894_o;
  wire _al_u897_o;
  wire _al_u898_o;
  wire _al_u899_o;
  wire _al_u900_o;
  wire _al_u903_o;
  wire _al_u904_o;
  wire _al_u906_o;
  wire _al_u908_o;
  wire _al_u909_o;
  wire _al_u912_o;
  wire _al_u913_o;
  wire _al_u914_o;
  wire _al_u916_o;
  wire _al_u920_o;
  wire _al_u922_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u926_o;
  wire _al_u927_o;
  wire _al_u930_o;
  wire _al_u931_o;
  wire _al_u932_o;
  wire _al_u933_o;
  wire _al_u935_o;
  wire _al_u938_o;
  wire _al_u939_o;
  wire _al_u940_o;
  wire _al_u941_o;
  wire _al_u942_o;
  wire _al_u944_o;
  wire _al_u945_o;
  wire _al_u946_o;
  wire _al_u948_o;
  wire _al_u951_o;
  wire _al_u952_o;
  wire _al_u953_o;
  wire _al_u954_o;
  wire _al_u955_o;
  wire _al_u956_o;
  wire _al_u958_o;
  wire _al_u960_o;
  wire _al_u963_o;
  wire _al_u964_o;
  wire _al_u965_o;
  wire _al_u966_o;
  wire _al_u967_o;
  wire _al_u968_o;
  wire _al_u970_o;
  wire _al_u972_o;
  wire _al_u975_o;
  wire _al_u976_o;
  wire _al_u977_o;
  wire _al_u978_o;
  wire _al_u979_o;
  wire _al_u980_o;
  wire _al_u982_o;
  wire _al_u984_o;
  wire _al_u987_o;
  wire _al_u988_o;
  wire _al_u989_o;
  wire _al_u990_o;
  wire _al_u991_o;
  wire _al_u992_o;
  wire _al_u994_o;
  wire _al_u996_o;
  wire _al_u999_o;
  wire \u1/c1 ;
  wire \u1/c11 ;
  wire \u1/c13 ;
  wire \u1/c3 ;
  wire \u1/c5 ;
  wire \u1/c7 ;
  wire \u1/c9 ;
  wire \u2/c1 ;
  wire \u2/c11 ;
  wire \u2/c13 ;
  wire \u2/c3 ;
  wire \u2/c5 ;
  wire \u2/c7 ;
  wire \u2/c9 ;
  wire \u_M0clkpll/clk0_buf ;  // al_ip/M0clkpll.v(34)
  wire \u_cmsdk_mcu/HWRITE ;  // ../RTL/cmsdk_mcu.v(106)
  wire \u_cmsdk_mcu/LOCKUPRESET ;  // ../RTL/cmsdk_mcu.v(86)
  wire \u_cmsdk_mcu/SYSRESETREQ ;  // ../RTL/cmsdk_mcu.v(78)
  wire \u_cmsdk_mcu/dbg_swdo ;  // ../RTL/cmsdk_mcu.v(166)
  wire \u_cmsdk_mcu/dbg_swdo_en ;  // ../RTL/cmsdk_mcu.v(165)
  wire \u_cmsdk_mcu/flash_hsel ;  // ../RTL/cmsdk_mcu.v(111)
  wire \u_cmsdk_mcu/n1 ;
  wire \u_cmsdk_mcu/sram_hsel ;  // ../RTL/cmsdk_mcu.v(117)
  wire \u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ;
  wire \u_cmsdk_mcu/u_ahb_ram/n16 ;
  wire \u_cmsdk_mcu/u_ahb_ram/we ;  // ../RTL/AHB2MEM.v(29)
  wire \u_cmsdk_mcu/u_ahb_rom/n16 ;
  wire \u_cmsdk_mcu/u_ahb_rom/we ;  // ../RTL/AHB2MEM.v(29)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ;  // ../RTL/cmsdk_mcu_clkctrl.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/nxt_hrst ;  // ../RTL/cmsdk_mcu_clkctrl.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ;  // ../RTL/cmsdk_mcu_clkctrl.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED ;  // ../RTL/cmsdk_mcu_system.v(171)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv ;  // ../RTL/cmsdk_mcu_system.v(80)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ;  // ../RTL/cmsdk_mcu_system.v(121)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hreadyout ;  // ../RTL/cmsdk_mcu_system.v(251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hsel ;  // ../RTL/cmsdk_mcu_system.v(250)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq ;  // ../RTL/cmsdk_mcu_system.v(342)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_hsel ;  // ../RTL/cmsdk_mcu_system.v(255)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/gpio1_hsel ;  // ../RTL/cmsdk_mcu_system.v(260)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/remap_ctrl ;  // ../RTL/cmsdk_mcu_system.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/sysctrl_hsel ;  // ../RTL/cmsdk_mcu_system.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel ;  // ../RTL/cmsdk_mcu_system.v(286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL ;  // ../RTL/cmsdk_ahb_gpio.v(75)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ;  // ../RTL/cmsdk_ahb_gpio.v(79)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ;  // ../RTL/cmsdk_ahb_gpio.v(77)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n101 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n103 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n105 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n107 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n109 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n111 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n113 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n115 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n117 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n119 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n121 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n123 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n125 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n127 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n129 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n144 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n146 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n148 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n150 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n152 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n154 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n156 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n158 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n160 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n162 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n164 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n166 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n168 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n170 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n172 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n174 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n189 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n191 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n193 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n195 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n197 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n199 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n201 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n203 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n205 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n207 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n209 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n211 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n213 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n215 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n217 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n219 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n234 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n236 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n238 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n240 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n242 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n244 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n246 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n248 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n250 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n252 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n254 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n256 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n258 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n260 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n262 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n264 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n271 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n273 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n275 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n277 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n279 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n281 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n283 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n285 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n287 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n289 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n291 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n293 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n295 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n297 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n299 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n301 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n54 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n56 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n58 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n60 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n62 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n64 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n66 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n68 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n70 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n72 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n74 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n76 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n78 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n80 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n82 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n84 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n99 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] ;  // ../RTL/cmsdk_ahb_gpio.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL ;  // ../RTL/cmsdk_ahb_gpio.v(75)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n101 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n103 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n105 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n107 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n109 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n111 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n113 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n115 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n117 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n119 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n121 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n123 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n125 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n127 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n129 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n144 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n146 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n148 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n150 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n152 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n154 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n156 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n158 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n160 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n162 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n164 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n166 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n168 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n170 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n172 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n174 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n189 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n191 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n193 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n195 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n197 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n199 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n201 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n203 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n205 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n207 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n209 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n211 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n213 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n215 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n217 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n219 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n234 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n236 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n238 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n240 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n242 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n244 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n246 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n248 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n250 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n252 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n254 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n256 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n258 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n260 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n262 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n264 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n271 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n273 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n275 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n277 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n279 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n281 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n283 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n285 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n287 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n289 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n291 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n293 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n295 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n297 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n299 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n301 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n54 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n56 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n58 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n60 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n62 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n64 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n66 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n68 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n70 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n72 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n74 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n76 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n78 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n80 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n82 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n84 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n99 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(266)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ;  // ../RTL/cmsdk_iop_gpio.v(514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ;  // ../RTL/cmsdk_iop_gpio.v(515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(105)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ;  // ../RTL/gpio.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n12_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ;  // ../RTL/cmsdk_apb_uart.v(76)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ;  // ../RTL/cmsdk_apb_uart.v(128)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b6_sel_is_13_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n106 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n114 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n117 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n31 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n40_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n46 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n48 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n50 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_txd ;  // ../RTL/cmsdk_apb_uart.v(163)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ;  // ../RTL/cmsdk_apb_uart.v(102)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun ;  // ../RTL/cmsdk_apb_uart.v(135)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ;  // ../RTL/cmsdk_apb_uart.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ;  // ../RTL/cmsdk_apb_uart.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full ;  // ../RTL/cmsdk_apb_uart.v(184)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun ;  // ../RTL/cmsdk_apb_uart.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ;  // ../RTL/cmsdk_apb_uart.v(172)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ;  // ../RTL/cmsdk_apb_uart.v(181)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ;  // ../RTL/cmsdk_apb_uart.v(177)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ;  // ../RTL/cmsdk_apb_uart.v(186)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1 ;  // ../RTL/cmsdk_apb_uart.v(168)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2 ;  // ../RTL/cmsdk_apb_uart.v(169)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ;  // ../RTL/cmsdk_apb_uart.v(161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun ;  // ../RTL/cmsdk_apb_uart.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ;  // ../RTL/cmsdk_apb_uart.v(154)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ;  // ../RTL/cmsdk_apb_uart.v(153)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_reg_txd ;  // ../RTL/cmsdk_apb_uart.v(164)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ;  // ../RTL/cmsdk_apb_uart.v(180)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ;  // ../RTL/cmsdk_apb_uart.v(103)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ;  // ../RTL/cmsdk_apb_uart.v(104)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ;  // ../RTL/cmsdk_apb_uart.v(106)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ;  // ../RTL/cmsdk_apb_uart.v(107)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ;  // ../RTL/cmsdk_apb_uart.v(108)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ;  // ../RTL/cmsdk_ahb_to_apb.v(88)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint ;  // ../RTL/cmsdk_apb_subsystem_m0ds.v(248)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ;  // ../RTL/cmsdk_mcu_sysctrl.v(116)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b6_sel_is_13_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_write ;  // ../RTL/cmsdk_mcu_sysctrl.v(280)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable ;  // ../RTL/cmsdk_mcu_sysctrl.v(121)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_write ;  // ../RTL/cmsdk_mcu_sysctrl.v(240)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ;  // ../RTL/cmsdk_mcu_sysctrl.v(309)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ;  // ../RTL/cmsdk_mcu_sysctrl.v(297)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable ;  // ../RTL/cmsdk_mcu_sysctrl.v(122)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED ;  // ../RTL/CORTEXM0INTEGRATION.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1047)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0mow6 ;  // ../RTL/cortexm0ds_logic.v(1141)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ;  // ../RTL/cortexm0ds_logic.v(371)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2cpw6 ;  // ../RTL/cortexm0ds_logic.v(1489)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ;  // ../RTL/cortexm0ds_logic.v(652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3biu6 ;  // ../RTL/cortexm0ds_logic.v(452)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ;  // ../RTL/cortexm0ds_logic.v(545)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4pow6 ;  // ../RTL/cortexm0ds_logic.v(1182)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A59pw6 ;  // ../RTL/cortexm0ds_logic.v(1450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(855)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1211)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ;  // ../RTL/cortexm0ds_logic.v(548)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad8pw6 ;  // ../RTL/cortexm0ds_logic.v(1440)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ;  // ../RTL/cortexm0ds_logic.v(602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(309)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 ;  // ../RTL/cortexm0ds_logic.v(376)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ;  // ../RTL/cortexm0ds_logic.v(283)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(738)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ai2ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(818)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aj1ju6 ;  // ../RTL/cortexm0ds_logic.v(805)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ;  // ../RTL/cortexm0ds_logic.v(524)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Akuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1255)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(860)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(392)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 ;  // ../RTL/cortexm0ds_logic.v(948)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ;  // ../RTL/cortexm0ds_logic.v(1229)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anciu6 ;  // ../RTL/cortexm0ds_logic.v(472)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(446)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ;  // ../RTL/cortexm0ds_logic.v(540)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqniu6 ;  // ../RTL/cortexm0ds_logic.v(621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ;  // ../RTL/cortexm0ds_logic.v(569)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Av3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ;  // ../RTL/cortexm0ds_logic.v(743)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awwow6 ;  // ../RTL/cortexm0ds_logic.v(1286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 ;  // ../RTL/cortexm0ds_logic.v(597)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ;  // ../RTL/cortexm0ds_logic.v(450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 ;  // ../RTL/cortexm0ds_logic.v(1007)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0iiu6 ;  // ../RTL/cortexm0ds_logic.v(544)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ;  // ../RTL/cortexm0ds_logic.v(424)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ;  // ../RTL/cortexm0ds_logic.v(1048)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4mow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1142)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6dow6 ;  // ../RTL/cortexm0ds_logic.v(1022)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8bow6 ;  // ../RTL/cortexm0ds_logic.v(996)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B91ju6 ;  // ../RTL/cortexm0ds_logic.v(801)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bagow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1064)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ;  // ../RTL/cortexm0ds_logic.v(601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 ;  // ../RTL/cortexm0ds_logic.v(588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bddow6 ;  // ../RTL/cortexm0ds_logic.v(1025)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 ;  // ../RTL/cortexm0ds_logic.v(736)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bg9iu6 ;  // ../RTL/cortexm0ds_logic.v(430)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(523)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 ;  // ../RTL/cortexm0ds_logic.v(710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ;  // ../RTL/cortexm0ds_logic.v(310)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bimow6 ;  // ../RTL/cortexm0ds_logic.v(1147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ;  // ../RTL/cortexm0ds_logic.v(684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bofiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(513)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ;  // ../RTL/cortexm0ds_logic.v(606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 ;  // ../RTL/cortexm0ds_logic.v(593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4pw6 ;  // ../RTL/cortexm0ds_logic.v(1392)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu2pw6 ;  // ../RTL/cortexm0ds_logic.v(1366)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwliu6 ;  // ../RTL/cortexm0ds_logic.v(596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxeow6 ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ;  // ../RTL/cortexm0ds_logic.v(851)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ;  // ../RTL/cortexm0ds_logic.v(1692)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 ;  // ../RTL/cortexm0ds_logic.v(1515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4iiu6 ;  // ../RTL/cortexm0ds_logic.v(546)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ;  // ../RTL/cortexm0ds_logic.v(345)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ;  // ../RTL/cortexm0ds_logic.v(600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 ;  // ../RTL/cortexm0ds_logic.v(1050)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8liu6 ;  // ../RTL/cortexm0ds_logic.v(587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C96pw6 ;  // ../RTL/cortexm0ds_logic.v(1411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ;  // ../RTL/cortexm0ds_logic.v(280)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(455)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchiu6 ;  // ../RTL/cortexm0ds_logic.v(535)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cemiu6 ;  // ../RTL/cortexm0ds_logic.v(603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cenow6 ;  // ../RTL/cortexm0ds_logic.v(1159)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ;  // ../RTL/cortexm0ds_logic.v(590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(858)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chkhu6 ;  // ../RTL/cortexm0ds_logic.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ciqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjiow6 ;  // ../RTL/cortexm0ds_logic.v(1094)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ;  // ../RTL/cortexm0ds_logic.v(325)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(780)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ;  // ../RTL/cortexm0ds_logic.v(949)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6 ;  // ../RTL/cortexm0ds_logic.v(1717)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqoiu6 ;  // ../RTL/cortexm0ds_logic.v(634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 ;  // ../RTL/cortexm0ds_logic.v(621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs7ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(889)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 ;  // ../RTL/cortexm0ds_logic.v(1164)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctliu6 ;  // ../RTL/cortexm0ds_logic.v(595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ;  // ../RTL/cortexm0ds_logic.v(475)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ;  // ../RTL/cortexm0ds_logic.v(556)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ;  // ../RTL/cortexm0ds_logic.v(891)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D14pw6 ;  // ../RTL/cortexm0ds_logic.v(1382)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ;  // ../RTL/cortexm0ds_logic.v(799)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ;  // ../RTL/cortexm0ds_logic.v(425)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ;  // ../RTL/cortexm0ds_logic.v(492)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(573)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1223)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ;  // ../RTL/cortexm0ds_logic.v(547)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(521)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbmiu6 ;  // ../RTL/cortexm0ds_logic.v(602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ;  // ../RTL/cortexm0ds_logic.v(776)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 ;  // ../RTL/cortexm0ds_logic.v(945)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ;  // ../RTL/cortexm0ds_logic.v(362)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgapw6 ;  // ../RTL/cortexm0ds_logic.v(1467)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ;  // ../RTL/cortexm0ds_logic.v(323)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ;  // ../RTL/cortexm0ds_logic.v(511)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6pw6 ;  // ../RTL/cortexm0ds_logic.v(1415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ;  // ../RTL/cortexm0ds_logic.v(947)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkeow6 ;  // ../RTL/cortexm0ds_logic.v(1041)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 ;  // ../RTL/cortexm0ds_logic.v(578)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ;  // ../RTL/cortexm0ds_logic.v(552)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ;  // ../RTL/cortexm0ds_logic.v(1202)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dooow6 ;  // ../RTL/cortexm0ds_logic.v(1176)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqfhu6 ;  // ../RTL/cortexm0ds_logic.v(125)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 ;  // ../RTL/cortexm0ds_logic.v(950)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ;  // ../RTL/cortexm0ds_logic.v(581)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drzow6 ;  // ../RTL/cortexm0ds_logic.v(1324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt4iu6 ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ;  // ../RTL/cortexm0ds_logic.v(1111)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ;  // ../RTL/cortexm0ds_logic.v(435)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzdow6 ;  // ../RTL/cortexm0ds_logic.v(1033)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ;  // ../RTL/cortexm0ds_logic.v(1610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(879)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ;  // ../RTL/cortexm0ds_logic.v(598)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2liu6 ;  // ../RTL/cortexm0ds_logic.v(585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ;  // ../RTL/cortexm0ds_logic.v(278)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yow6 ;  // ../RTL/cortexm0ds_logic.v(1303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5jow6 ;  // ../RTL/cortexm0ds_logic.v(1102)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8miu6 ;  // ../RTL/cortexm0ds_logic.v(601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9mow6 ;  // ../RTL/cortexm0ds_logic.v(1144)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ea7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(944)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 ;  // ../RTL/cortexm0ds_logic.v(668)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eazow6 ;  // ../RTL/cortexm0ds_logic.v(1318)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ;  // ../RTL/cortexm0ds_logic.v(1011)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eciiu6 ;  // ../RTL/cortexm0ds_logic.v(549)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1466)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(523)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef7ju6 ;  // ../RTL/cortexm0ds_logic.v(884)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ;  // ../RTL/cortexm0ds_logic.v(390)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eidow6 ;  // ../RTL/cortexm0ds_logic.v(1027)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejaju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(926)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ;  // ../RTL/cortexm0ds_logic.v(1482)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejcow6 ;  // ../RTL/cortexm0ds_logic.v(1014)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ekhiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(538)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ;  // ../RTL/cortexm0ds_logic.v(1594)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emmiu6 ;  // ../RTL/cortexm0ds_logic.v(606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(767)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epciu6 ;  // ../RTL/cortexm0ds_logic.v(473)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 ;  // ../RTL/cortexm0ds_logic.v(567)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ;  // ../RTL/cortexm0ds_logic.v(286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eq4pw6 ;  // ../RTL/cortexm0ds_logic.v(1391)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ;  // ../RTL/cortexm0ds_logic.v(1204)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eriow6 ;  // ../RTL/cortexm0ds_logic.v(1097)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(421)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eukhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 ;  // ../RTL/cortexm0ds_logic.v(582)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(569)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1219)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 ;  // ../RTL/cortexm0ds_logic.v(811)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ;  // ../RTL/cortexm0ds_logic.v(1034)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ;  // ../RTL/cortexm0ds_logic.v(664)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F15pw6 ;  // ../RTL/cortexm0ds_logic.v(1395)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 ;  // ../RTL/cortexm0ds_logic.v(1690)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F42iu6 ;  // ../RTL/cortexm0ds_logic.v(332)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(880)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ;  // ../RTL/cortexm0ds_logic.v(412)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ;  // ../RTL/cortexm0ds_logic.v(1249)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ;  // ../RTL/cortexm0ds_logic.v(774)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7zhu6 ;  // ../RTL/cortexm0ds_logic.v(293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ;  // ../RTL/cortexm0ds_logic.v(373)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 ;  // ../RTL/cortexm0ds_logic.v(1210)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faoiu6 ;  // ../RTL/cortexm0ds_logic.v(628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fdfow6 ;  // ../RTL/cortexm0ds_logic.v(1052)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ;  // ../RTL/cortexm0ds_logic.v(657)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1213)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 ;  // ../RTL/cortexm0ds_logic.v(282)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ;  // ../RTL/cortexm0ds_logic.v(644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ;  // ../RTL/cortexm0ds_logic.v(631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkliu6 ;  // ../RTL/cortexm0ds_logic.v(592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ;  // ../RTL/cortexm0ds_logic.v(1602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fllow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1135)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(935)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ;  // ../RTL/cortexm0ds_logic.v(1594)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ;  // ../RTL/cortexm0ds_logic.v(646)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ;  // ../RTL/cortexm0ds_logic.v(740)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(989)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(781)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 ;  // ../RTL/cortexm0ds_logic.v(394)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ;  // ../RTL/cortexm0ds_logic.v(488)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fucow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1018)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fviow6 ;  // ../RTL/cortexm0ds_logic.v(1099)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx9ow6 ;  // ../RTL/cortexm0ds_logic.v(979)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fy8ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(966)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ;  // ../RTL/cortexm0ds_logic.v(597)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ;  // ../RTL/cortexm0ds_logic.v(584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0phu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0pow6 ;  // ../RTL/cortexm0ds_logic.v(1181)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 ;  // ../RTL/cortexm0ds_logic.v(981)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2miu6 ;  // ../RTL/cortexm0ds_logic.v(598)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 ;  // ../RTL/cortexm0ds_logic.v(492)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 ;  // ../RTL/cortexm0ds_logic.v(1009)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xow6 ;  // ../RTL/cortexm0ds_logic.v(1290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7aiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(440)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ;  // ../RTL/cortexm0ds_logic.v(801)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 ;  // ../RTL/cortexm0ds_logic.v(1077)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(507)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc6ow6 ;  // ../RTL/cortexm0ds_logic.v(931)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gcjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(562)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd4pw6 ;  // ../RTL/cortexm0ds_logic.v(1386)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdjow6 ;  // ../RTL/cortexm0ds_logic.v(1105)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ;  // ../RTL/cortexm0ds_logic.v(1199)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(999)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 ;  // ../RTL/cortexm0ds_logic.v(804)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gggow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1066)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gglhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(832)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ;  // ../RTL/cortexm0ds_logic.v(364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4pw6 ;  // ../RTL/cortexm0ds_logic.v(1389)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ;  // ../RTL/cortexm0ds_logic.v(1014)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ;  // ../RTL/cortexm0ds_logic.v(1202)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 ;  // ../RTL/cortexm0ds_logic.v(739)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ;  // ../RTL/cortexm0ds_logic.v(445)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(312)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpeow6 ;  // ../RTL/cortexm0ds_logic.v(1043)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1230)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 ;  // ../RTL/cortexm0ds_logic.v(767)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1217)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwhhu6 ;  // ../RTL/cortexm0ds_logic.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwkiu6 ;  // ../RTL/cortexm0ds_logic.v(583)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gy3ju6 ;  // ../RTL/cortexm0ds_logic.v(838)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ;  // ../RTL/cortexm0ds_logic.v(1625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00pw6 ;  // ../RTL/cortexm0ds_logic.v(1328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1zhu6 ;  // ../RTL/cortexm0ds_logic.v(290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3bpw6 ;  // ../RTL/cortexm0ds_logic.v(1476)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(829)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha4pw6 ;  // ../RTL/cortexm0ds_logic.v(1385)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ;  // ../RTL/cortexm0ds_logic.v(454)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 ;  // ../RTL/cortexm0ds_logic.v(1653)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 ;  // ../RTL/cortexm0ds_logic.v(998)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbpow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1185)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(522)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcuiu6 ;  // ../RTL/cortexm0ds_logic.v(709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1146)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 ;  // ../RTL/cortexm0ds_logic.v(1068)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ;  // ../RTL/cortexm0ds_logic.v(592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(948)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hndow6 ;  // ../RTL/cortexm0ds_logic.v(1029)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoiiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(553)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(540)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ;  // ../RTL/cortexm0ds_logic.v(964)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ;  // ../RTL/cortexm0ds_logic.v(595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ;  // ../RTL/cortexm0ds_logic.v(769)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1018)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ;  // ../RTL/cortexm0ds_logic.v(556)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(449)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(543)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hy1pw6 ;  // ../RTL/cortexm0ds_logic.v(1354)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ;  // ../RTL/cortexm0ds_logic.v(610)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ;  // ../RTL/cortexm0ds_logic.v(316)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0pw6 ;  // ../RTL/cortexm0ds_logic.v(1341)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hzliu6 ;  // ../RTL/cortexm0ds_logic.v(597)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 ;  // ../RTL/cortexm0ds_logic.v(731)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ;  // ../RTL/cortexm0ds_logic.v(893)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(786)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I46ju6 ;  // ../RTL/cortexm0ds_logic.v(867)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ;  // ../RTL/cortexm0ds_logic.v(492)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ;  // ../RTL/cortexm0ds_logic.v(854)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ;  // ../RTL/cortexm0ds_logic.v(1674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1210)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(279)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7cow6 ;  // ../RTL/cortexm0ds_logic.v(1010)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ;  // ../RTL/cortexm0ds_logic.v(815)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ;  // ../RTL/cortexm0ds_logic.v(1653)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I98ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(895)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia0ju6 ;  // ../RTL/cortexm0ds_logic.v(789)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 ;  // ../RTL/cortexm0ds_logic.v(588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ;  // ../RTL/cortexm0ds_logic.v(1599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 ;  // ../RTL/cortexm0ds_logic.v(682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ;  // ../RTL/cortexm0ds_logic.v(575)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ;  // ../RTL/cortexm0ds_logic.v(843)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idkow6 ;  // ../RTL/cortexm0ds_logic.v(1119)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 ;  // ../RTL/cortexm0ds_logic.v(1599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iecow6 ;  // ../RTL/cortexm0ds_logic.v(1012)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iexow6 ;  // ../RTL/cortexm0ds_logic.v(1293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/If3pw6 ;  // ../RTL/cortexm0ds_logic.v(1374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ;  // ../RTL/cortexm0ds_logic.v(591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ;  // ../RTL/cortexm0ds_logic.v(1147)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ;  // ../RTL/cortexm0ds_logic.v(1612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ;  // ../RTL/cortexm0ds_logic.v(739)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ;  // ../RTL/cortexm0ds_logic.v(820)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inniu6 ;  // ../RTL/cortexm0ds_logic.v(620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Io9ow6 ;  // ../RTL/cortexm0ds_logic.v(976)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipliu6 ;  // ../RTL/cortexm0ds_logic.v(594)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqriu6 ;  // ../RTL/cortexm0ds_logic.v(674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1231)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ;  // ../RTL/cortexm0ds_logic.v(937)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isbpw6 ;  // ../RTL/cortexm0ds_logic.v(1485)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/It3iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(354)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itbow6 ;  // ../RTL/cortexm0ds_logic.v(1004)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ;  // ../RTL/cortexm0ds_logic.v(529)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivmiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1246)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(397)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 ;  // ../RTL/cortexm0ds_logic.v(1515)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3row6 ;  // ../RTL/cortexm0ds_logic.v(1209)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(746)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(826)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5pow6 ;  // ../RTL/cortexm0ds_logic.v(1183)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(319)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J77ju6 ;  // ../RTL/cortexm0ds_logic.v(881)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 ;  // ../RTL/cortexm0ds_logic.v(1674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ;  // ../RTL/cortexm0ds_logic.v(494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1050)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8ziu6 ;  // ../RTL/cortexm0ds_logic.v(774)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9eow6 ;  // ../RTL/cortexm0ds_logic.v(1037)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(574)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 ;  // ../RTL/cortexm0ds_logic.v(293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ;  // ../RTL/cortexm0ds_logic.v(374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jajiu6 ;  // ../RTL/cortexm0ds_logic.v(561)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 ;  // ../RTL/cortexm0ds_logic.v(655)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(829)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ;  // ../RTL/cortexm0ds_logic.v(1105)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jc3pw6 ;  // ../RTL/cortexm0ds_logic.v(1372)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ;  // ../RTL/cortexm0ds_logic.v(1185)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ;  // ../RTL/cortexm0ds_logic.v(871)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 ;  // ../RTL/cortexm0ds_logic.v(1146)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgeow6 ;  // ../RTL/cortexm0ds_logic.v(1040)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ;  // ../RTL/cortexm0ds_logic.v(1612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhyow6 ;  // ../RTL/cortexm0ds_logic.v(1307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ;  // ../RTL/cortexm0ds_logic.v(631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjwow6 ;  // ../RTL/cortexm0ds_logic.v(1281)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkhow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1081)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ;  // ../RTL/cortexm0ds_logic.v(605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(847)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ;  // ../RTL/cortexm0ds_logic.v(353)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jr1ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(808)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvow6 ;  // ../RTL/cortexm0ds_logic.v(1271)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ;  // ../RTL/cortexm0ds_logic.v(1615)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvdow6 ;  // ../RTL/cortexm0ds_logic.v(1032)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ;  // ../RTL/cortexm0ds_logic.v(1609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxow6 ;  // ../RTL/cortexm0ds_logic.v(1300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 ;  // ../RTL/cortexm0ds_logic.v(449)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6 ;  // ../RTL/cortexm0ds_logic.v(1645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy2pw6 ;  // ../RTL/cortexm0ds_logic.v(1367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy9iu6 ;  // ../RTL/cortexm0ds_logic.v(436)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzmiu6 ;  // ../RTL/cortexm0ds_logic.v(611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ;  // ../RTL/cortexm0ds_logic.v(745)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 ;  // ../RTL/cortexm0ds_logic.v(1007)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ;  // ../RTL/cortexm0ds_logic.v(425)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ;  // ../RTL/cortexm0ds_logic.v(612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(968)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ;  // ../RTL/cortexm0ds_logic.v(386)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(373)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1210)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8iiu6 ;  // ../RTL/cortexm0ds_logic.v(547)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ;  // ../RTL/cortexm0ds_logic.v(896)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kb9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(971)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ;  // ../RTL/cortexm0ds_logic.v(870)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kctow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 ;  // ../RTL/cortexm0ds_logic.v(630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kikhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 ;  // ../RTL/cortexm0ds_logic.v(578)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 ;  // ../RTL/cortexm0ds_logic.v(672)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(846)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ;  // ../RTL/cortexm0ds_logic.v(1028)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 ;  // ../RTL/cortexm0ds_logic.v(552)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ;  // ../RTL/cortexm0ds_logic.v(1202)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kp1pw6 ;  // ../RTL/cortexm0ds_logic.v(1351)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq0pw6 ;  // ../RTL/cortexm0ds_logic.v(1338)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ;  // ../RTL/cortexm0ds_logic.v(407)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krkiu6 ;  // ../RTL/cortexm0ds_logic.v(581)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kt4iu6 ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktwiu6 ;  // ../RTL/cortexm0ds_logic.v(742)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 ;  // ../RTL/cortexm0ds_logic.v(1005)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1192)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kv9iu6 ;  // ../RTL/cortexm0ds_logic.v(435)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ;  // ../RTL/cortexm0ds_logic.v(516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1260)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(784)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzkhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0how6 ;  // ../RTL/cortexm0ds_logic.v(1074)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ;  // ../RTL/cortexm0ds_logic.v(611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vow6 ;  // ../RTL/cortexm0ds_logic.v(1261)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ;  // ../RTL/cortexm0ds_logic.v(1613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L27pw6 ;  // ../RTL/cortexm0ds_logic.v(1422)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L3sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(372)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ;  // ../RTL/cortexm0ds_logic.v(1653)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1251)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9mow6 ;  // ../RTL/cortexm0ds_logic.v(1144)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 ;  // ../RTL/cortexm0ds_logic.v(1674)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ;  // ../RTL/cortexm0ds_logic.v(668)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ;  // ../RTL/cortexm0ds_logic.v(281)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ;  // ../RTL/cortexm0ds_logic.v(1199)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1092)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf1iu6 ;  // ../RTL/cortexm0ds_logic.v(322)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1066)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(484)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(832)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1482)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ;  // ../RTL/cortexm0ds_logic.v(551)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ll2pw6 ;  // ../RTL/cortexm0ds_logic.v(1362)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(988)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ;  // ../RTL/cortexm0ds_logic.v(325)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 ;  // ../RTL/cortexm0ds_logic.v(1717)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ;  // ../RTL/cortexm0ds_logic.v(1680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0pw6 ;  // ../RTL/cortexm0ds_logic.v(1336)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 ;  // ../RTL/cortexm0ds_logic.v(580)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 ;  // ../RTL/cortexm0ds_logic.v(1136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqcow6 ;  // ../RTL/cortexm0ds_logic.v(1017)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 ;  // ../RTL/cortexm0ds_logic.v(541)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 ;  // ../RTL/cortexm0ds_logic.v(809)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls9pw6 ;  // ../RTL/cortexm0ds_logic.v(1459)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ;  // ../RTL/cortexm0ds_logic.v(315)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 ;  // ../RTL/cortexm0ds_logic.v(952)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ;  // ../RTL/cortexm0ds_logic.v(824)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ;  // ../RTL/cortexm0ds_logic.v(1034)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M14ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ;  // ../RTL/cortexm0ds_logic.v(371)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 ;  // ../RTL/cortexm0ds_logic.v(745)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2cow6 ;  // ../RTL/cortexm0ds_logic.v(1008)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ;  // ../RTL/cortexm0ds_logic.v(574)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ;  // ../RTL/cortexm0ds_logic.v(293)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1211)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(828)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1078)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdfow6 ;  // ../RTL/cortexm0ds_logic.v(1052)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ;  // ../RTL/cortexm0ds_logic.v(563)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(831)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(899)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mj8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ;  // ../RTL/cortexm0ds_logic.v(1068)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmiu6 ;  // ../RTL/cortexm0ds_logic.v(605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjnow6 ;  // ../RTL/cortexm0ds_logic.v(1161)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjtiu6 ;  // ../RTL/cortexm0ds_logic.v(698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(873)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ml6pw6 ;  // ../RTL/cortexm0ds_logic.v(1416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 ;  // ../RTL/cortexm0ds_logic.v(1510)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(566)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 ;  // ../RTL/cortexm0ds_logic.v(659)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 ;  // ../RTL/cortexm0ds_logic.v(285)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ;  // ../RTL/cortexm0ds_logic.v(1593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpgiu6 ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ;  // ../RTL/cortexm0ds_logic.v(620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mq1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrfow6 ;  // ../RTL/cortexm0ds_logic.v(1057)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ;  // ../RTL/cortexm0ds_logic.v(1689)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt6ow6 ;  // ../RTL/cortexm0ds_logic.v(938)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mtrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1218)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ;  // ../RTL/cortexm0ds_logic.v(316)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ;  // ../RTL/cortexm0ds_logic.v(397)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzkiu6 ;  // ../RTL/cortexm0ds_logic.v(584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0phu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(892)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ;  // ../RTL/cortexm0ds_logic.v(773)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N45ju6 ;  // ../RTL/cortexm0ds_logic.v(853)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ;  // ../RTL/cortexm0ds_logic.v(1183)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(481)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(575)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(562)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3ju6 ;  // ../RTL/cortexm0ds_logic.v(830)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 ;  // ../RTL/cortexm0ds_logic.v(604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhlhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(565)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(926)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkxow6 ;  // ../RTL/cortexm0ds_logic.v(1295)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nn8iu6 ;  // ../RTL/cortexm0ds_logic.v(419)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(949)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npghu6 ;  // ../RTL/cortexm0ds_logic.v(127)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(848)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(448)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 ;  // ../RTL/cortexm0ds_logic.v(715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ;  // ../RTL/cortexm0ds_logic.v(1689)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ;  // ../RTL/cortexm0ds_logic.v(978)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 ;  // ../RTL/cortexm0ds_logic.v(396)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 ;  // ../RTL/cortexm0ds_logic.v(1046)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1220)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nycow6 ;  // ../RTL/cortexm0ds_logic.v(1020)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxow6 ;  // ../RTL/cortexm0ds_logic.v(1300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 ;  // ../RTL/cortexm0ds_logic.v(825)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O16iu6 ;  // ../RTL/cortexm0ds_logic.v(384)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ;  // ../RTL/cortexm0ds_logic.v(371)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4bow6 ;  // ../RTL/cortexm0ds_logic.v(995)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(426)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ;  // ../RTL/cortexm0ds_logic.v(361)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oaxow6 ;  // ../RTL/cortexm0ds_logic.v(1292)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(998)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocniu6 ;  // ../RTL/cortexm0ds_logic.v(616)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(509)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ;  // ../RTL/cortexm0ds_logic.v(1065)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oe7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1240)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Of5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(857)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogdow6 ;  // ../RTL/cortexm0ds_logic.v(1026)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogqiu6 ;  // ../RTL/cortexm0ds_logic.v(657)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ;  // ../RTL/cortexm0ds_logic.v(831)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ;  // ../RTL/cortexm0ds_logic.v(363)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6 ;  // ../RTL/cortexm0ds_logic.v(1706)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok7ju6 ;  // ../RTL/cortexm0ds_logic.v(886)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 ;  // ../RTL/cortexm0ds_logic.v(951)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(837)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 ;  // ../RTL/cortexm0ds_logic.v(649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ;  // ../RTL/cortexm0ds_logic.v(636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhhu6 ;  // ../RTL/cortexm0ds_logic.v(129)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhow6 ;  // ../RTL/cortexm0ds_logic.v(1086)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oy8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ;  // ../RTL/cortexm0ds_logic.v(451)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ;  // ../RTL/cortexm0ds_logic.v(1007)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ;  // ../RTL/cortexm0ds_logic.v(344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ;  // ../RTL/cortexm0ds_logic.v(1625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P22iu6 ;  // ../RTL/cortexm0ds_logic.v(331)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1249)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 ;  // ../RTL/cortexm0ds_logic.v(586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ;  // ../RTL/cortexm0ds_logic.v(828)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(453)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8aiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(440)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 ;  // ../RTL/cortexm0ds_logic.v(721)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P92iu6 ;  // ../RTL/cortexm0ds_logic.v(334)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 ;  // ../RTL/cortexm0ds_logic.v(614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pa7ju6 ;  // ../RTL/cortexm0ds_logic.v(882)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pagow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1064)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ;  // ../RTL/cortexm0ds_logic.v(575)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ;  // ../RTL/cortexm0ds_logic.v(1676)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyow6 ;  // ../RTL/cortexm0ds_logic.v(1306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peqow6 ;  // ../RTL/cortexm0ds_logic.v(1199)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 ;  // ../RTL/cortexm0ds_logic.v(1612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 ;  // ../RTL/cortexm0ds_logic.v(323)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(417)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1254)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ;  // ../RTL/cortexm0ds_logic.v(778)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pj7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(947)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ;  // ../RTL/cortexm0ds_logic.v(765)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ;  // ../RTL/cortexm0ds_logic.v(846)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ;  // ../RTL/cortexm0ds_logic.v(1028)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ;  // ../RTL/cortexm0ds_logic.v(1717)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 ;  // ../RTL/cortexm0ds_logic.v(365)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmoiu6 ;  // ../RTL/cortexm0ds_logic.v(633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ;  // ../RTL/cortexm0ds_logic.v(406)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1231)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Prdow6 ;  // ../RTL/cortexm0ds_logic.v(1030)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ;  // ../RTL/cortexm0ds_logic.v(542)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(809)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwfow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1059)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxlow6 ;  // ../RTL/cortexm0ds_logic.v(1140)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 ;  // ../RTL/cortexm0ds_logic.v(677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(570)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(289)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q07ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(879)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1fow6 ;  // ../RTL/cortexm0ds_logic.v(1048)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ;  // ../RTL/cortexm0ds_logic.v(1035)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 ;  // ../RTL/cortexm0ds_logic.v(1712)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(840)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ;  // ../RTL/cortexm0ds_logic.v(652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5hiu6 ;  // ../RTL/cortexm0ds_logic.v(533)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 ;  // ../RTL/cortexm0ds_logic.v(600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7uow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1250)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1237)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ;  // ../RTL/cortexm0ds_logic.v(1619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ;  // ../RTL/cortexm0ds_logic.v(374)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(468)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ;  // ../RTL/cortexm0ds_logic.v(655)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(829)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1373)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ;  // ../RTL/cortexm0ds_logic.v(1689)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 ;  // ../RTL/cortexm0ds_logic.v(442)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1079)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qgkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj2ju6 ;  // ../RTL/cortexm0ds_logic.v(819)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(899)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1456)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ;  // ../RTL/cortexm0ds_logic.v(418)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ;  // ../RTL/cortexm0ds_logic.v(1707)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qodow6 ;  // ../RTL/cortexm0ds_logic.v(1029)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qoyow6 ;  // ../RTL/cortexm0ds_logic.v(1310)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ;  // ../RTL/cortexm0ds_logic.v(541)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ;  // ../RTL/cortexm0ds_logic.v(528)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1058)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ;  // ../RTL/cortexm0ds_logic.v(1045)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxbow6 ;  // ../RTL/cortexm0ds_logic.v(1006)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ;  // ../RTL/cortexm0ds_logic.v(637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qy2pw6 ;  // ../RTL/cortexm0ds_logic.v(1367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ;  // ../RTL/cortexm0ds_logic.v(798)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ;  // ../RTL/cortexm0ds_logic.v(838)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0ghu6 ;  // ../RTL/cortexm0ds_logic.v(125)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ;  // ../RTL/cortexm0ds_logic.v(519)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1075)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R47ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(880)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5eiu6 ;  // ../RTL/cortexm0ds_logic.v(493)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(828)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ;  // ../RTL/cortexm0ds_logic.v(441)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9wow6 ;  // ../RTL/cortexm0ds_logic.v(1278)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ;  // ../RTL/cortexm0ds_logic.v(1676)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rb7ju6 ;  // ../RTL/cortexm0ds_logic.v(883)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ;  // ../RTL/cortexm0ds_logic.v(589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ;  // ../RTL/cortexm0ds_logic.v(776)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1213)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ;  // ../RTL/cortexm0ds_logic.v(524)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(617)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhoow6 ;  // ../RTL/cortexm0ds_logic.v(1174)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ;  // ../RTL/cortexm0ds_logic.v(604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1241)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ;  // ../RTL/cortexm0ds_logic.v(779)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk5ju6 ;  // ../RTL/cortexm0ds_logic.v(859)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ;  // ../RTL/cortexm0ds_logic.v(1651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ;  // ../RTL/cortexm0ds_logic.v(578)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1228)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ;  // ../RTL/cortexm0ds_logic.v(298)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ;  // ../RTL/cortexm0ds_logic.v(1483)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 ;  // ../RTL/cortexm0ds_logic.v(552)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro1ju6 ;  // ../RTL/cortexm0ds_logic.v(807)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro2pw6 ;  // ../RTL/cortexm0ds_logic.v(1364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 ;  // ../RTL/cortexm0ds_logic.v(1618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs5pw6 ;  // ../RTL/cortexm0ds_logic.v(1405)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(287)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rt4pw6 ;  // ../RTL/cortexm0ds_logic.v(1392)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 ;  // ../RTL/cortexm0ds_logic.v(823)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1192)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvniu6 ;  // ../RTL/cortexm0ds_logic.v(623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw8iu6 ;  // ../RTL/cortexm0ds_logic.v(422)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwgow6 ;  // ../RTL/cortexm0ds_logic.v(1072)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ;  // ../RTL/cortexm0ds_logic.v(1643)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(477)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S02iu6 ;  // ../RTL/cortexm0ds_logic.v(330)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1tiu6 ;  // ../RTL/cortexm0ds_logic.v(692)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(772)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 ;  // ../RTL/cortexm0ds_logic.v(572)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S63iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(346)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6ihu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ow6 ;  // ../RTL/cortexm0ds_logic.v(957)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ;  // ../RTL/cortexm0ds_logic.v(1212)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 ;  // ../RTL/cortexm0ds_logic.v(281)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ;  // ../RTL/cortexm0ds_logic.v(455)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdoiu6 ;  // ../RTL/cortexm0ds_logic.v(629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdwow6 ;  // ../RTL/cortexm0ds_logic.v(1279)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ;  // ../RTL/cortexm0ds_logic.v(323)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh7ow6 ;  // ../RTL/cortexm0ds_logic.v(947)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjkhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ;  // ../RTL/cortexm0ds_logic.v(1201)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smnow6 ;  // ../RTL/cortexm0ds_logic.v(1162)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 ;  // ../RTL/cortexm0ds_logic.v(406)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ;  // ../RTL/cortexm0ds_logic.v(580)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Spyhu6 ;  // ../RTL/cortexm0ds_logic.v(286)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ;  // ../RTL/cortexm0ds_logic.v(835)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ;  // ../RTL/cortexm0ds_logic.v(1004)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ;  // ../RTL/cortexm0ds_logic.v(1618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1259)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 ;  // ../RTL/cortexm0ds_logic.v(1650)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 ;  // ../RTL/cortexm0ds_logic.v(289)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ;  // ../RTL/cortexm0ds_logic.v(824)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6 ;  // ../RTL/cortexm0ds_logic.v(1625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ;  // ../RTL/cortexm0ds_logic.v(852)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 ;  // ../RTL/cortexm0ds_logic.v(290)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zow6 ;  // ../RTL/cortexm0ds_logic.v(1315)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T14ju6 ;  // ../RTL/cortexm0ds_logic.v(839)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(826)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ;  // ../RTL/cortexm0ds_logic.v(800)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ;  // ../RTL/cortexm0ds_logic.v(1592)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ;  // ../RTL/cortexm0ds_logic.v(1676)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6ziu6 ;  // ../RTL/cortexm0ds_logic.v(774)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ;  // ../RTL/cortexm0ds_logic.v(854)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 ;  // ../RTL/cortexm0ds_logic.v(1198)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ;  // ../RTL/cortexm0ds_logic.v(415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 ;  // ../RTL/cortexm0ds_logic.v(295)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ;  // ../RTL/cortexm0ds_logic.v(1716)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tj1iu6 ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ;  // ../RTL/cortexm0ds_logic.v(1707)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkfow6 ;  // ../RTL/cortexm0ds_logic.v(1055)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tktow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ;  // ../RTL/cortexm0ds_logic.v(1706)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 ;  // ../RTL/cortexm0ds_logic.v(659)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 ;  // ../RTL/cortexm0ds_logic.v(1216)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(821)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 ;  // ../RTL/cortexm0ds_logic.v(1605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsriu6 ;  // ../RTL/cortexm0ds_logic.v(675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 ;  // ../RTL/cortexm0ds_logic.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttmhu6 ;  // ../RTL/cortexm0ds_logic.v(143)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1018)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tw2iu6 ;  // ../RTL/cortexm0ds_logic.v(342)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ;  // ../RTL/cortexm0ds_logic.v(423)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ;  // ../RTL/cortexm0ds_logic.v(490)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1234)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ;  // ../RTL/cortexm0ds_logic.v(344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0oiu6 ;  // ../RTL/cortexm0ds_logic.v(625)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ;  // ../RTL/cortexm0ds_logic.v(424)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 ;  // ../RTL/cortexm0ds_logic.v(705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U28iu6 ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ;  // ../RTL/cortexm0ds_logic.v(279)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 ;  // ../RTL/cortexm0ds_logic.v(734)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U73iu6 ;  // ../RTL/cortexm0ds_logic.v(346)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 ;  // ../RTL/cortexm0ds_logic.v(708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ;  // ../RTL/cortexm0ds_logic.v(414)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U99ow6 ;  // ../RTL/cortexm0ds_logic.v(970)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ;  // ../RTL/cortexm0ds_logic.v(843)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ;  // ../RTL/cortexm0ds_logic.v(362)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 ;  // ../RTL/cortexm0ds_logic.v(1467)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uehiu6 ;  // ../RTL/cortexm0ds_logic.v(536)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uf9iu6 ;  // ../RTL/cortexm0ds_logic.v(430)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufkhu6 ;  // ../RTL/cortexm0ds_logic.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(417)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ugmiu6 ;  // ../RTL/cortexm0ds_logic.v(604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ;  // ../RTL/cortexm0ds_logic.v(1678)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4ju6 ;  // ../RTL/cortexm0ds_logic.v(846)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ;  // ../RTL/cortexm0ds_logic.v(565)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1483)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ;  // ../RTL/cortexm0ds_logic.v(1652)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ;  // ../RTL/cortexm0ds_logic.v(619)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 ;  // ../RTL/cortexm0ds_logic.v(713)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ;  // ../RTL/cortexm0ds_logic.v(593)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 ;  // ../RTL/cortexm0ds_logic.v(687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ;  // ../RTL/cortexm0ds_logic.v(1687)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1230)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqyow6 ;  // ../RTL/cortexm0ds_logic.v(1311)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ;  // ../RTL/cortexm0ds_logic.v(367)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ;  // ../RTL/cortexm0ds_logic.v(822)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(448)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utgiu6 ;  // ../RTL/cortexm0ds_logic.v(528)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu8iu6 ;  // ../RTL/cortexm0ds_logic.v(422)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(978)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 ;  // ../RTL/cortexm0ds_logic.v(596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ;  // ../RTL/cortexm0ds_logic.v(690)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwdpw6 ;  // ../RTL/cortexm0ds_logic.v(1514)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzow6 ;  // ../RTL/cortexm0ds_logic.v(1327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux5iu6 ;  // ../RTL/cortexm0ds_logic.v(383)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1488)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ;  // ../RTL/cortexm0ds_logic.v(557)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ;  // ../RTL/cortexm0ds_logic.v(450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V17ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(941)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1low6 ;  // ../RTL/cortexm0ds_logic.v(1128)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1221)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1115)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 ;  // ../RTL/cortexm0ds_logic.v(358)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3cow6 ;  // ../RTL/cortexm0ds_logic.v(1008)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ;  // ../RTL/cortexm0ds_logic.v(265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V4phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52iu6 ;  // ../RTL/cortexm0ds_logic.v(332)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ;  // ../RTL/cortexm0ds_logic.v(426)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5oow6 ;  // ../RTL/cortexm0ds_logic.v(1169)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V77pw6 ;  // ../RTL/cortexm0ds_logic.v(1424)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ;  // ../RTL/cortexm0ds_logic.v(1011)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1091)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 ;  // ../RTL/cortexm0ds_logic.v(603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 ;  // ../RTL/cortexm0ds_logic.v(777)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ;  // ../RTL/cortexm0ds_logic.v(577)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(538)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(618)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(834)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(460)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ;  // ../RTL/cortexm0ds_logic.v(1203)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ;  // ../RTL/cortexm0ds_logic.v(740)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voxow6 ;  // ../RTL/cortexm0ds_logic.v(1297)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 ;  // ../RTL/cortexm0ds_logic.v(1709)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 ;  // ../RTL/cortexm0ds_logic.v(1589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 ;  // ../RTL/cortexm0ds_logic.v(634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 ;  // ../RTL/cortexm0ds_logic.v(1715)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ;  // ../RTL/cortexm0ds_logic.v(1606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 ;  // ../RTL/cortexm0ds_logic.v(314)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs7pw6 ;  // ../RTL/cortexm0ds_logic.v(1432)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 ;  // ../RTL/cortexm0ds_logic.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vu5iu6 ;  // ../RTL/cortexm0ds_logic.v(382)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ;  // ../RTL/cortexm0ds_logic.v(475)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ;  // ../RTL/cortexm0ds_logic.v(556)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vwapw6 ;  // ../RTL/cortexm0ds_logic.v(1474)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ;  // ../RTL/cortexm0ds_logic.v(436)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ;  // ../RTL/cortexm0ds_logic.v(1645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1167)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ;  // ../RTL/cortexm0ds_logic.v(1588)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ;  // ../RTL/cortexm0ds_logic.v(344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1wow6 ;  // ../RTL/cortexm0ds_logic.v(1275)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W38pw6 ;  // ../RTL/cortexm0ds_logic.v(1436)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ;  // ../RTL/cortexm0ds_logic.v(305)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W48ow6 ;  // ../RTL/cortexm0ds_logic.v(955)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 ;  // ../RTL/cortexm0ds_logic.v(1517)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 ;  // ../RTL/cortexm0ds_logic.v(1049)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 ;  // ../RTL/cortexm0ds_logic.v(680)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 ;  // ../RTL/cortexm0ds_logic.v(1584)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 ;  // ../RTL/cortexm0ds_logic.v(453)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ;  // ../RTL/cortexm0ds_logic.v(1010)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9lhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ;  // ../RTL/cortexm0ds_logic.v(789)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 ;  // ../RTL/cortexm0ds_logic.v(1711)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 ;  // ../RTL/cortexm0ds_logic.v(602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ;  // ../RTL/cortexm0ds_logic.v(308)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbkhu6 ;  // ../RTL/cortexm0ds_logic.v(136)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(856)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ;  // ../RTL/cortexm0ds_logic.v(456)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ;  // ../RTL/cortexm0ds_logic.v(1702)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfihu6 ;  // ../RTL/cortexm0ds_logic.v(131)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 ;  // ../RTL/cortexm0ds_logic.v(724)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ;  // ../RTL/cortexm0ds_logic.v(791)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(973)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 ;  // ../RTL/cortexm0ds_logic.v(1067)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 ;  // ../RTL/cortexm0ds_logic.v(1638)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ;  // ../RTL/cortexm0ds_logic.v(765)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wk5pw6 ;  // ../RTL/cortexm0ds_logic.v(1402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkciu6 ;  // ../RTL/cortexm0ds_logic.v(472)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ;  // ../RTL/cortexm0ds_logic.v(565)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ;  // ../RTL/cortexm0ds_logic.v(1015)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlxow6 ;  // ../RTL/cortexm0ds_logic.v(1296)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 ;  // ../RTL/cortexm0ds_logic.v(726)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Womiu6 ;  // ../RTL/cortexm0ds_logic.v(607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ;  // ../RTL/cortexm0ds_logic.v(300)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr6ow6 ;  // ../RTL/cortexm0ds_logic.v(937)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrcpw6 ;  // ../RTL/cortexm0ds_logic.v(1499)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(368)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtbow6 ;  // ../RTL/cortexm0ds_logic.v(1005)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 ;  // ../RTL/cortexm0ds_logic.v(729)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv8pw6 ;  // ../RTL/cortexm0ds_logic.v(1447)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv9ow6 ;  // ../RTL/cortexm0ds_logic.v(979)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ;  // ../RTL/cortexm0ds_logic.v(1645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ww6ju6 ;  // ../RTL/cortexm0ds_logic.v(877)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1140)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ;  // ../RTL/cortexm0ds_logic.v(771)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wy4ju6 ;  // ../RTL/cortexm0ds_logic.v(851)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wydow6 ;  // ../RTL/cortexm0ds_logic.v(1033)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyhhu6 ;  // ../RTL/cortexm0ds_logic.v(130)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ;  // ../RTL/cortexm0ds_logic.v(1649)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 ;  // ../RTL/cortexm0ds_logic.v(664)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ;  // ../RTL/cortexm0ds_logic.v(370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 ;  // ../RTL/cortexm0ds_logic.v(651)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ;  // ../RTL/cortexm0ds_logic.v(504)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ;  // ../RTL/cortexm0ds_logic.v(585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2zhu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(291)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 ;  // ../RTL/cortexm0ds_logic.v(1621)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X53pw6 ;  // ../RTL/cortexm0ds_logic.v(1370)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 ;  // ../RTL/cortexm0ds_logic.v(158)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ;  // ../RTL/cortexm0ds_logic.v(1606)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X62pw6 ;  // ../RTL/cortexm0ds_logic.v(1357)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ;  // ../RTL/cortexm0ds_logic.v(613)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X71pw6 ;  // ../RTL/cortexm0ds_logic.v(1344)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ;  // ../RTL/cortexm0ds_logic.v(1697)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 ;  // ../RTL/cortexm0ds_logic.v(600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ;  // ../RTL/cortexm0ds_logic.v(1614)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80pw6 ;  // ../RTL/cortexm0ds_logic.v(1331)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87iu6 ;  // ../RTL/cortexm0ds_logic.v(400)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87pw6 ;  // ../RTL/cortexm0ds_logic.v(1425)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(842)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 ;  // ../RTL/cortexm0ds_logic.v(1714)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1011)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbiiu6 ;  // ../RTL/cortexm0ds_logic.v(548)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(816)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ;  // ../RTL/cortexm0ds_logic.v(1630)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 ;  // ../RTL/cortexm0ds_logic.v(1636)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 ;  // ../RTL/cortexm0ds_logic.v(1705)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ;  // ../RTL/cortexm0ds_logic.v(1603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ;  // ../RTL/cortexm0ds_logic.v(1628)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfliu6 ;  // ../RTL/cortexm0ds_logic.v(590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ;  // ../RTL/cortexm0ds_logic.v(390)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ;  // ../RTL/cortexm0ds_logic.v(364)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 ;  // ../RTL/cortexm0ds_logic.v(925)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ;  // ../RTL/cortexm0ds_logic.v(457)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ;  // ../RTL/cortexm0ds_logic.v(1585)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ;  // ../RTL/cortexm0ds_logic.v(645)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(325)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ;  // ../RTL/cortexm0ds_logic.v(1627)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xneow6 ;  // ../RTL/cortexm0ds_logic.v(1042)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ;  // ../RTL/cortexm0ds_logic.v(1682)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ;  // ../RTL/cortexm0ds_logic.v(1640)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ;  // ../RTL/cortexm0ds_logic.v(1204)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ;  // ../RTL/cortexm0ds_logic.v(1684)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1378)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqpow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1191)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ;  // ../RTL/cortexm0ds_logic.v(528)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ;  // ../RTL/cortexm0ds_logic.v(1675)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ;  // ../RTL/cortexm0ds_logic.v(327)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ;  // ../RTL/cortexm0ds_logic.v(608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1245)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 ;  // ../RTL/cortexm0ds_logic.v(1622)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(769)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ;  // ../RTL/cortexm0ds_logic.v(301)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ;  // ../RTL/cortexm0ds_logic.v(938)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 ;  // ../RTL/cortexm0ds_logic.v(1695)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 ;  // ../RTL/cortexm0ds_logic.v(1633)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6 ;  // ../RTL/cortexm0ds_logic.v(1691)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ;  // ../RTL/cortexm0ds_logic.v(450)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 ;  // ../RTL/cortexm0ds_logic.v(1600)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ;  // ../RTL/cortexm0ds_logic.v(1608)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xyohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xz9ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(980)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ;  // ../RTL/cortexm0ds_logic.v(1167)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ;  // ../RTL/cortexm0ds_logic.v(1708)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ;  // ../RTL/cortexm0ds_logic.v(558)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ;  // ../RTL/cortexm0ds_logic.v(1195)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xow6 ;  // ../RTL/cortexm0ds_logic.v(1288)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 ;  // ../RTL/cortexm0ds_logic.v(1641)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2hiu6 ;  // ../RTL/cortexm0ds_logic.v(532)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2phu6 ;  // ../RTL/cortexm0ds_logic.v(157)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y32pw6 ;  // ../RTL/cortexm0ds_logic.v(1356)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3niu6 ;  // ../RTL/cortexm0ds_logic.v(612)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ;  // ../RTL/cortexm0ds_logic.v(787)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y41pw6 ;  // ../RTL/cortexm0ds_logic.v(1343)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 ;  // ../RTL/cortexm0ds_logic.v(599)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ;  // ../RTL/cortexm0ds_logic.v(306)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50pw6 ;  // ../RTL/cortexm0ds_logic.v(1330)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 ;  // ../RTL/cortexm0ds_logic.v(1637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 ;  // ../RTL/cortexm0ds_logic.v(138)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 ;  // ../RTL/cortexm0ds_logic.v(586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 ;  // ../RTL/cortexm0ds_logic.v(1683)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7cpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1491)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7yow6 ;  // ../RTL/cortexm0ds_logic.v(1304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ;  // ../RTL/cortexm0ds_logic.v(360)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ;  // ../RTL/cortexm0ds_logic.v(1590)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 ;  // ../RTL/cortexm0ds_logic.v(1685)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ;  // ../RTL/cortexm0ds_logic.v(347)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(802)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 ;  // ../RTL/cortexm0ds_logic.v(1265)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ;  // ../RTL/cortexm0ds_logic.v(415)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc0pw6 ;  // ../RTL/cortexm0ds_logic.v(1333)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ;  // ../RTL/cortexm0ds_logic.v(402)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ;  // ../RTL/cortexm0ds_logic.v(589)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1239)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yd7ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(945)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ;  // ../RTL/cortexm0ds_logic.v(576)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1494)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ;  // ../RTL/cortexm0ds_logic.v(1620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ;  // ../RTL/cortexm0ds_logic.v(1013)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfiiu6 ;  // ../RTL/cortexm0ds_logic.v(550)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 ;  // ../RTL/cortexm0ds_logic.v(1200)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yg3iu6 ;  // ../RTL/cortexm0ds_logic.v(350)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yh8ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(898)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(324)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(885)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(417)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yj8ow6 ;  // ../RTL/cortexm0ds_logic.v(961)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 ;  // ../RTL/cortexm0ds_logic.v(1632)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjtow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1242)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykkiu6 ;  // ../RTL/cortexm0ds_logic.v(579)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1229)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ;  // ../RTL/cortexm0ds_logic.v(566)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ;  // ../RTL/cortexm0ds_logic.v(1624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ;  // ../RTL/cortexm0ds_logic.v(365)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 ;  // ../RTL/cortexm0ds_logic.v(740)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6 ;  // ../RTL/cortexm0ds_logic.v(1611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(352)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynwow6 ;  // ../RTL/cortexm0ds_logic.v(1283)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ;  // ../RTL/cortexm0ds_logic.v(807)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 ;  // ../RTL/cortexm0ds_logic.v(1644)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(527)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 ;  // ../RTL/cortexm0ds_logic.v(137)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ;  // ../RTL/cortexm0ds_logic.v(620)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ;  // ../RTL/cortexm0ds_logic.v(781)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ;  // ../RTL/cortexm0ds_logic.v(1677)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ;  // ../RTL/cortexm0ds_logic.v(849)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysihu6 ;  // ../RTL/cortexm0ds_logic.v(132)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ;  // ../RTL/cortexm0ds_logic.v(836)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ;  // ../RTL/cortexm0ds_logic.v(1688)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ;  // ../RTL/cortexm0ds_logic.v(1700)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yuiow6 ;  // ../RTL/cortexm0ds_logic.v(1099)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ;  // ../RTL/cortexm0ds_logic.v(810)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv9pw6 ;  // ../RTL/cortexm0ds_logic.v(1460)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ;  // ../RTL/cortexm0ds_logic.v(1699)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ;  // ../RTL/cortexm0ds_logic.v(529)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ;  // ../RTL/cortexm0ds_logic.v(1587)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ;  // ../RTL/cortexm0ds_logic.v(329)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ;  // ../RTL/cortexm0ds_logic.v(1686)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 ;  // ../RTL/cortexm0ds_logic.v(1639)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ;  // ../RTL/cortexm0ds_logic.v(1602)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yy7ow6 ;  // ../RTL/cortexm0ds_logic.v(953)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ;  // ../RTL/cortexm0ds_logic.v(1635)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 ;  // ../RTL/cortexm0ds_logic.v(303)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 ;  // ../RTL/cortexm0ds_logic.v(664)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 ;  // ../RTL/cortexm0ds_logic.v(1601)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ;  // ../RTL/cortexm0ds_logic.v(1604)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z08ju6_lutinv ;  // ../RTL/cortexm0ds_logic.v(892)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0niu6 ;  // ../RTL/cortexm0ds_logic.v(611)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(411)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18pw6 ;  // ../RTL/cortexm0ds_logic.v(1435)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ;  // ../RTL/cortexm0ds_logic.v(505)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 ;  // ../RTL/cortexm0ds_logic.v(598)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 ;  // ../RTL/cortexm0ds_logic.v(304)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ;  // ../RTL/cortexm0ds_logic.v(1631)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 ;  // ../RTL/cortexm0ds_logic.v(1516)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2fow6 ;  // ../RTL/cortexm0ds_logic.v(1048)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(941)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3sow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1222)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z4kow6 ;  // ../RTL/cortexm0ds_logic.v(1116)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 ;  // ../RTL/cortexm0ds_logic.v(359)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 ;  // ../RTL/cortexm0ds_logic.v(1626)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6iow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1090)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ;  // ../RTL/cortexm0ds_logic.v(1681)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ;  // ../RTL/cortexm0ds_logic.v(1623)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ;  // ../RTL/cortexm0ds_logic.v(1586)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ;  // ../RTL/cortexm0ds_logic.v(307)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ;  // ../RTL/cortexm0ds_logic.v(1698)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ;  // ../RTL/cortexm0ds_logic.v(1596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Za6pw6 ;  // ../RTL/cortexm0ds_logic.v(1412)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 ;  // ../RTL/cortexm0ds_logic.v(562)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zccow6 ;  // ../RTL/cortexm0ds_logic.v(1012)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 ;  // ../RTL/cortexm0ds_logic.v(1701)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 ;  // ../RTL/cortexm0ds_logic.v(1647)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ;  // ../RTL/cortexm0ds_logic.v(1605)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 ;  // ../RTL/cortexm0ds_logic.v(139)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ;  // ../RTL/cortexm0ds_logic.v(884)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8iu6 ;  // ../RTL/cortexm0ds_logic.v(416)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfgow6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1066)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 ;  // ../RTL/cortexm0ds_logic.v(603)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ;  // ../RTL/cortexm0ds_logic.v(403)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ;  // ../RTL/cortexm0ds_logic.v(1634)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ;  // ../RTL/cortexm0ds_logic.v(1642)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(778)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zi5iu6 ;  // ../RTL/cortexm0ds_logic.v(377)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 ;  // ../RTL/cortexm0ds_logic.v(1696)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 ;  // ../RTL/cortexm0ds_logic.v(1704)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zokiu6 ;  // ../RTL/cortexm0ds_logic.v(580)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zpkow6 ;  // ../RTL/cortexm0ds_logic.v(1123)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ;  // ../RTL/cortexm0ds_logic.v(1648)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(541)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ;  // ../RTL/cortexm0ds_logic.v(1591)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 ;  // ../RTL/cortexm0ds_logic.v(1679)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ;  // ../RTL/cortexm0ds_logic.v(328)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ;  // ../RTL/cortexm0ds_logic.v(609)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ;  // ../RTL/cortexm0ds_logic.v(1607)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ;  // ../RTL/cortexm0ds_logic.v(596)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 ;  // ../RTL/cortexm0ds_logic.v(1710)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 ;  // ../RTL/cortexm0ds_logic.v(583)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ;  // ../RTL/cortexm0ds_logic.v(302)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ;  // ../RTL/cortexm0ds_logic.v(1500)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ;  // ../RTL/cortexm0ds_logic.v(1595)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ;  // ../RTL/cortexm0ds_logic.v(1629)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ;  // ../RTL/cortexm0ds_logic.v(1703)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 ;  // ../RTL/cortexm0ds_logic.v(637)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ;  // ../RTL/cortexm0ds_logic.v(624)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzohu6 ;  // ../RTL/cortexm0ds_logic.v(156)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c31 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[12]_i1[12]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[16]_i1[16]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[1]_i1[1]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[21]_i1[21]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[27]_i1[27]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[3]_i1[3]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[5]_i1[5]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[12]_i1[12]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[15]_i1[15]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[1]_i1[1]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[5]_i1[5]_o_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_14 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_16 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_17 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_18 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_20 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_21 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_22 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_24 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_25 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_26 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_27 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_28 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_29 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_30 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_31 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_0 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_10 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_12 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_13 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_2 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_4 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_6 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_8 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_9 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n267 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3436 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n590 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c11 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c15 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c19 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c23 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c1 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c3 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c5 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c7 ;
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ;  // ../RTL/cortexm0ds_logic.v(70)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ;  // ../RTL/cortexm0ds_logic.v(117)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ;  // ../RTL/cortexm0ds_logic.v(71)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] ;  // ../RTL/cortexm0ds_logic.v(67)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ;  // ../RTL/cortexm0ds_logic.v(69)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ;  // ../RTL/cortexm0ds_logic.v(118)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] ;  // ../RTL/cortexm0ds_logic.v(68)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] ;  // ../RTL/cortexm0ds_logic.v(53)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] ;  // ../RTL/cortexm0ds_logic.v(63)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ;  // ../RTL/cortexm0ds_logic.v(64)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] ;  // ../RTL/cortexm0ds_logic.v(65)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] ;  // ../RTL/cortexm0ds_logic.v(66)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] ;  // ../RTL/cortexm0ds_logic.v(54)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] ;  // ../RTL/cortexm0ds_logic.v(55)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] ;  // ../RTL/cortexm0ds_logic.v(56)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] ;  // ../RTL/cortexm0ds_logic.v(57)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] ;  // ../RTL/cortexm0ds_logic.v(58)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] ;  // ../RTL/cortexm0ds_logic.v(59)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] ;  // ../RTL/cortexm0ds_logic.v(60)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] ;  // ../RTL/cortexm0ds_logic.v(61)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] ;  // ../RTL/cortexm0ds_logic.v(62)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ;  // ../RTL/cortexm0ds_logic.v(116)
  wire \u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ;  // ../RTL/cmsdk_ahb_cs_rom_table.v(157)
  wire uart0_txd_pad;  // ../RTL/M0demo.v(20)
  wire uart0_txen_pad;  // ../RTL/M0demo.v(21)

  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u100 (
    .do({open_n1,open_n2,open_n3,\u_cmsdk_mcu/p0_out [10]}),
    .ts(\u_cmsdk_mcu/p0_outen [10]),
    .opad(P0[10]));  // ../RTL/cmsdk_mcu_pin_mux.v(136)
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    //.LUT1("(~D*~(~A*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000001111),
    .INIT_LUT1(16'b0000000011101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1000|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b2  (
    .a({_al_u996_o,open_n16}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [2],open_n17}),
    .c({_al_u999_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [2]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,b_pad_gpio_porta_pad[2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1000_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [2]}),
    .q({open_n34,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [2]}));  // ../RTL/gpio_ctrl.v(184)
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*~A*~(C*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*~A*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1001|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b2  (
    .a({_al_u1000_o,open_n35}),
    .b({_al_u945_o,open_n36}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [2],_al_u2490_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/HWDATA [2]}),
    .mi({open_n40,\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1001_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n193 }),
    .q({open_n55,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [2]}));  // ../RTL/gpio_apbif.v(383)
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011111111110101),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011111111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1002|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2],open_n56}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [2],open_n57}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2492_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [2]}),
    .mi({open_n61,\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n148 }),
    .q({open_n76,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [2]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1003|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2],open_n77}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [2],open_n78}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2496_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [2]}),
    .mi({open_n89,\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1003_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n58 }),
    .q({open_n93,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2]}));  // ../RTL/gpio_apbif.v(323)
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1004|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b2  (
    .b({_al_u1002_o,_al_u1004_o}),
    .c({_al_u1003_o,_al_u1006_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u566_o,_al_u1001_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1004_o,open_n108}),
    .q({open_n112,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [2]}));  // ../RTL/gpio_apbif.v(453)
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTF1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTG1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000001110111),
    .INIT_LUTF1(16'b0000000010101100),
    .INIT_LUTG0(16'b0010000001110111),
    .INIT_LUTG1(16'b0000000010101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1005|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2],\u_cmsdk_mcu/HWDATA [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 }),
    .mi({open_n116,\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b2/B1_0 ,_al_u3342_o}),
    .q({open_n131,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]}));  // ../RTL/gpio_apbif.v(262)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B*A))"),
    //.LUTF1("(~D*~(~C*~B*A))"),
    //.LUTG0("(~D*~(~C*~B*A))"),
    //.LUTG1("(~D*~(~C*~B*A))"),
    .INIT_LUTF0(16'b0000000011111101),
    .INIT_LUTF1(16'b0000000011111101),
    .INIT_LUTG0(16'b0000000011111101),
    .INIT_LUTG1(16'b0000000011111101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1006|_al_u982  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b2/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b4/B1_0 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .f({_al_u1006_o,_al_u982_o}));
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~(C*B)))"),
    //.LUTF1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTG0("(A*~(D*~(C*B)))"),
    //.LUTG1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000010101010),
    .INIT_LUTF1(16'b1010100000001000),
    .INIT_LUTG0(16'b1000000010101010),
    .INIT_LUTG1(16'b1010100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1008|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b1  (
    .a({_al_u470_o,_al_u3456_o}),
    .b({b_pad_gpio_porta_pad[1],\u_cmsdk_mcu/HWDATA [1]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 }),
    .mi({open_n159,\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1008_o,_al_u3457_o}),
    .q({open_n174,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]}));  // ../RTL/gpio_apbif.v(262)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u101 (
    .do({open_n176,open_n177,open_n178,\u_cmsdk_mcu/p0_out [9]}),
    .ts(\u_cmsdk_mcu/p0_outen [9]),
    .opad(P0[9]));  // ../RTL/cmsdk_mcu_pin_mux.v(135)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(B*A)))"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(~C*~(D*~(B*A)))"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b0000100000001111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1010|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [1],\u_cmsdk_mcu/HWDATA [1]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [1],_al_u3075_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [1]}),
    .mi({open_n194,\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1010_o,_al_u3076_o}),
    .q({open_n209,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [1]}));  // ../RTL/gpio_apbif.v(323)
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000001111),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1011|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b1  (
    .a({_al_u1010_o,open_n210}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1],open_n211}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [1]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,b_pad_gpio_porta_pad[1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1011_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [1]}),
    .q({open_n228,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [1]}));  // ../RTL/gpio_ctrl.v(184)
  // ../RTL/gpio_apbif.v(343)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~A*~(C*~(~D*~B)))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~A*~(C*~(~D*~B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000010100010101),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1012|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b1  (
    .a({_al_u1008_o,open_n229}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [1],open_n230}),
    .c({_al_u1011_o,_al_u2496_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1],\u_cmsdk_mcu/HWDATA [1]}),
    .mi({open_n234,\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1012_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n56 }),
    .q({open_n249,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1]}));  // ../RTL/gpio_apbif.v(343)
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1013|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [1],open_n252}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,_al_u2492_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({_al_u945_o,\u_cmsdk_mcu/HWDATA [1]}),
    .mi({open_n256,\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1013_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n146 }),
    .q({open_n271,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [1]}));  // ../RTL/gpio_apbif.v(383)
  // ../RTL/gpio_apbif.v(242)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000010101100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000010101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1014|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1],open_n272}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1],open_n273}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2490_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [1]}),
    .mi({open_n277,\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b1/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n191 }),
    .q({open_n292,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1]}));  // ../RTL/gpio_apbif.v(242)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B*A))"),
    //.LUTF1("(~D*~(~C*~B*A))"),
    //.LUTG0("(~D*~(~C*~B*A))"),
    //.LUTG1("(~D*~(~C*~B*A))"),
    .INIT_LUTF0(16'b0000000011111101),
    .INIT_LUTF1(16'b0000000011111101),
    .INIT_LUTG0(16'b0000000011111101),
    .INIT_LUTG1(16'b0000000011111101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1015|_al_u970  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b1/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b5/B1_0 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .f({_al_u1015_o,_al_u970_o}));
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1016|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1],open_n317}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [1],open_n318}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2494_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [1]}),
    .mi({open_n329,\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1016_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n101 }),
    .q({open_n333,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [1]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1017|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [1],open_n334}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [1],open_n335}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,_al_u3076_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1017_o,open_n349}),
    .q({open_n353,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [1]}));  // ../RTL/gpio_ctrl.v(248)
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(~D*~A)))"),
    //.LUT1("(A*~(B*~(D*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000111),
    .INIT_LUT1(16'b1010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1018|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b1  (
    .a({_al_u1015_o,_al_u1012_o}),
    .b({_al_u566_o,_al_u1013_o}),
    .c({_al_u1016_o,_al_u1018_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u1017_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1018_o,open_n366}),
    .q({open_n370,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [1]}));  // ../RTL/gpio_apbif.v(453)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u102 (
    .do({open_n372,open_n373,open_n374,\u_cmsdk_mcu/p0_out [8]}),
    .ts(\u_cmsdk_mcu/p0_outen [8]),
    .opad(P0[8]));  // ../RTL/cmsdk_mcu_pin_mux.v(134)
  // ../RTL/gpio_apbif.v(242)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1010100000001000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1010100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1020|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b0  (
    .a({_al_u470_o,open_n387}),
    .b({b_pad_gpio_porta_pad[0],_al_u467_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0],_al_u472_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }),
    .mi({open_n391,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1020_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 }),
    .q({open_n406,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0]}));  // ../RTL/gpio_apbif.v(242)
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100100000001000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1022|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [0],open_n407}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0],_al_u692_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [0],_al_u467_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }),
    .mi({open_n411,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 }),
    .q({open_n426,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0]}));  // ../RTL/gpio_apbif.v(303)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~D*~C*~(~B*A))"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~D*~C*~(~B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000001101),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000000001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1023|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u692_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .mi({open_n430,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1023_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 }),
    .q({open_n445,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0]}));  // ../RTL/gpio_apbif.v(323)
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(D*~A*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1025|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b0  (
    .a({_al_u1024_o,open_n446}),
    .b({_al_u945_o,_al_u945_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }),
    .mi({open_n457,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1025_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 }),
    .q({open_n461,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }));  // ../RTL/gpio_apbif.v(383)
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0011111111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1026|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0],open_n462}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [0],_al_u692_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u1048_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }),
    .mi({open_n473,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1026_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 }),
    .q({open_n477,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [0]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_apbif.v(343)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1027|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0],open_n478}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [0],_al_u692_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u571_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }),
    .mi({open_n489,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1027_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 }),
    .q({open_n493,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [0]}));  // ../RTL/gpio_apbif.v(343)
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1028|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b0  (
    .b({_al_u1026_o,_al_u1028_o}),
    .c({_al_u1027_o,_al_u1030_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u566_o,_al_u1025_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1028_o,open_n508}),
    .q({open_n512,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [0]}));  // ../RTL/gpio_apbif.v(453)
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C@D)"),
    //.LUTF1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG0("~(C@D)"),
    //.LUTG1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000001111),
    .INIT_LUTF1(16'b0000000010101100),
    .INIT_LUTG0(16'b1111000000001111),
    .INIT_LUTG1(16'b0000000010101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1029|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0],open_n513}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0],open_n514}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [0]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,b_pad_gpio_porta_pad[0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b0/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [0]}),
    .q({open_n535,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [0]}));  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u103 (
    .do({open_n537,open_n538,open_n539,\u_cmsdk_mcu/p0_out [7]}),
    .ts(\u_cmsdk_mcu/p0_outen [7]),
    .opad(P0[7]));  // ../RTL/cmsdk_mcu_pin_mux.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B*A))"),
    //.LUT1("(~D*~(~C*~B*A))"),
    .INIT_LUT0(16'b0000000011111101),
    .INIT_LUT1(16'b0000000011111101),
    .MODE("LOGIC"))
    \_al_u1030|_al_u958  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b0/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b6/B1_0 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .f({_al_u1030_o,_al_u958_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(B*~(~D*C)))"),
    //.LUTF1("(D*~C*B*~A)"),
    //.LUTG0("~(A*~(B*~(~D*C)))"),
    //.LUTG1("(D*~C*B*~A)"),
    .INIT_LUTF0(16'b1101110101011101),
    .INIT_LUTF1(16'b0000010000000000),
    .INIT_LUTG0(16'b1101110101011101),
    .INIT_LUTG1(16'b0000010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1032|_al_u638  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ,_al_u637_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2],_al_u379_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv }),
    .f({_al_u1032_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~B*A)"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(D*C*~B*A)"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1033|_al_u636  (
    .a({open_n596,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full }),
    .f({_al_u1033_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(A*~(D*B)))"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b0000110100000101),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u1034|_al_u1039  (
    .a({open_n621,_al_u1034_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1],uart0_txen_pad}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full }),
    .f({_al_u1034_o,_al_u1039_o}));
  // ../RTL/cmsdk_apb_uart.v(445)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~D*~(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1035|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b2  (
    .b({_al_u1034_o,open_n644}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ),
    .clk(XTAL1_wire),
    .d({_al_u1033_o,_al_u1035_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1035_o,open_n657}),
    .q({open_n661,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]}));  // ../RTL/cmsdk_apb_uart.v(445)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u104 (
    .do({open_n663,open_n664,open_n665,\u_cmsdk_mcu/p0_out [6]}),
    .ts(\u_cmsdk_mcu/p0_outen [6]),
    .opad(P0[6]));  // ../RTL/cmsdk_mcu_pin_mux.v(132)
  // ../RTL/cmsdk_apb_uart.v(445)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b0001000100111111),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b0001000100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1040|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b0  (
    .a({_al_u1033_o,open_n678}),
    .b({_al_u1039_o,open_n679}),
    .c({_al_u1034_o,_al_u1040_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [0],_al_u1032_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1040_o,open_n696}),
    .q({open_n700,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]}));  // ../RTL/cmsdk_apb_uart.v(445)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*B*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1046|_al_u6830  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ,open_n703}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ,_al_u6830_o}));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u105 (
    .do({open_n729,open_n730,open_n731,\u_cmsdk_mcu/p0_out [5]}),
    .ts(\u_cmsdk_mcu/p0_outen [5]),
    .opad(P0[5]));  // ../RTL/cmsdk_mcu_pin_mux.v(131)
  // ../RTL/cortexm0ds_logic.v(18948)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~D*C*B*~A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~D*C*B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000000001000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1050|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lxwax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] }),
    .mi({open_n747,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ll2pw6 }),
    .q({open_n763,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] }));  // ../RTL/cortexm0ds_logic.v(18948)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*~A)"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(D*~C*B*~A)"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b0000010000000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000010000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1051|_al_u1880  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }));
  // ../RTL/cortexm0ds_logic.v(18922)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1053|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uhvax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] }),
    .mi({open_n798,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,_al_u1193_o}),
    .q({open_n803,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] }));  // ../RTL/cortexm0ds_logic.v(18922)
  // ../RTL/cortexm0ds_logic.v(17849)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1054|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkxpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] }),
    .mi({open_n814,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,_al_u1073_o}),
    .q({open_n819,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] }));  // ../RTL/cortexm0ds_logic.v(17849)
  // ../RTL/cortexm0ds_logic.v(18900)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1055|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bauax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] }),
    .mi({open_n830,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({_al_u1055_o,_al_u714_o}),
    .q({open_n835,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[0] }));  // ../RTL/cortexm0ds_logic.v(18900)
  // ../RTL/cortexm0ds_logic.v(18711)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~D*C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1056|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oykax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] }),
    .mi({open_n846,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,_al_u1058_o}),
    .q({open_n851,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] }));  // ../RTL/cortexm0ds_logic.v(18711)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~A)"),
    //.LUT1("(~D*C*~B*~A)"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000000000010000),
    .MODE("LOGIC"))
    \_al_u1057|_al_u1879  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*~A)"),
    //.LUT1("(~D*~C*B*A)"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"))
    \_al_u1059|_al_u1874  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u106 (
    .do({open_n893,open_n894,open_n895,\u_cmsdk_mcu/p0_out [4]}),
    .ts(\u_cmsdk_mcu/p0_outen [4]),
    .opad(P0[4]));  // ../RTL/cmsdk_mcu_pin_mux.v(130)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*~A)"),
    //.LUTF1("(~D*~C*B*~A)"),
    //.LUTG0("(D*C*B*~A)"),
    //.LUTG1("(~D*~C*B*~A)"),
    .INIT_LUTF0(16'b0100000000000000),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0100000000000000),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1060|_al_u1872  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }));
  // ../RTL/cortexm0ds_logic.v(18797)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1062|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kloax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X53pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .b({_al_u1055_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1058_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1061_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] }),
    .mi({open_n935,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ,_al_u1061_o}),
    .q({open_n951,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] }));  // ../RTL/cortexm0ds_logic.v(18797)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1063|_al_u5988  (
    .a({open_n952,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 }),
    .b({open_n953,_al_u607_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ,_al_u932_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [0],_al_u5988_o}));
  // ../RTL/cortexm0ds_logic.v(18820)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1066|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvpax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] }),
    .mi({open_n988,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u1066_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0pow6 }),
    .q({open_n993,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[2] }));  // ../RTL/cortexm0ds_logic.v(18820)
  // ../RTL/cortexm0ds_logic.v(18792)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1068|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mboax6_reg  (
    .a({_al_u1064_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({_al_u1065_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({_al_u1066_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu2pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] }),
    .mi({open_n997,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ,_al_u1065_o}),
    .q({open_n1013,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[2] }));  // ../RTL/cortexm0ds_logic.v(18792)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1069|_al_u872  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [3]}));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u107 (
    .do({open_n1043,open_n1044,open_n1045,\u_cmsdk_mcu/p0_out [3]}),
    .ts(\u_cmsdk_mcu/p0_outen [3]),
    .opad(P0[3]));  // ../RTL/cmsdk_mcu_pin_mux.v(129)
  // ../RTL/cortexm0ds_logic.v(18817)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1070|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eppax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] }),
    .mi({open_n1061,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({_al_u1070_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cenow6 }),
    .q({open_n1077,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[10] }));  // ../RTL/cortexm0ds_logic.v(18817)
  // ../RTL/cortexm0ds_logic.v(18845)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1074|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8rax6_reg  (
    .a({_al_u1070_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .b({_al_u1071_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ll2pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1073_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] }),
    .mi({open_n1081,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 ,_al_u1071_o}),
    .q({open_n1097,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[10] }));  // ../RTL/cortexm0ds_logic.v(18845)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1075|_al_u818  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [27]}));
  // ../RTL/cortexm0ds_logic.v(18974)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1076|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3yax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] }),
    .mi({open_n1129,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1076_o,_al_u870_o}),
    .q({open_n1145,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[3] }));  // ../RTL/cortexm0ds_logic.v(18974)
  // ../RTL/cortexm0ds_logic.v(18798)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1078|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jnoax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] }),
    .mi({open_n1149,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1078_o,_al_u868_o}),
    .q({open_n1165,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[3] }));  // ../RTL/cortexm0ds_logic.v(18798)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u108 (
    .do({open_n1167,open_n1168,open_n1169,\u_cmsdk_mcu/p0_out [2]}),
    .ts(\u_cmsdk_mcu/p0_outen [2]),
    .opad(P0[2]));  // ../RTL/cmsdk_mcu_pin_mux.v(128)
  // ../RTL/cortexm0ds_logic.v(17544)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1080|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktppw6_reg  (
    .a({_al_u1076_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({_al_u1077_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({_al_u1078_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1079_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] }),
    .mi({open_n1192,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ,_al_u1079_o}),
    .q({open_n1197,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[3] }));  // ../RTL/cortexm0ds_logic.v(17544)
  // ../RTL/cortexm0ds_logic.v(19776)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1082|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cm7bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,open_n1198}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,open_n1199}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv }),
    .mi({open_n1203,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .f({_al_u1082_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 }),
    .q({open_n1219,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] }));  // ../RTL/cortexm0ds_logic.v(19776)
  // ../RTL/cortexm0ds_logic.v(19768)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1083|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C67bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] }),
    .mi({open_n1230,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .f({_al_u1083_o,_al_u900_o}),
    .q({open_n1235,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[11] }));  // ../RTL/cortexm0ds_logic.v(19768)
  // ../RTL/cortexm0ds_logic.v(18928)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1084|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rtvax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] }),
    .mi({open_n1239,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y32pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X53pw6 }),
    .q({open_n1255,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[0] }));  // ../RTL/cortexm0ds_logic.v(18928)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u1086|_al_u1164  (
    .a({_al_u1082_o,_al_u1160_o}),
    .b({_al_u1083_o,_al_u1161_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y32pw6 ,_al_u1162_o}),
    .d({_al_u1085_o,_al_u1163_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 }));
  // ../RTL/cortexm0ds_logic.v(18821)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1088|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxpax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] }),
    .mi({open_n1286,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1088_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4pow6 }),
    .q({open_n1291,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[4] }));  // ../RTL/cortexm0ds_logic.v(18821)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u109 (
    .do({open_n1293,open_n1294,open_n1295,\u_cmsdk_mcu/p0_out [1]}),
    .ts(\u_cmsdk_mcu/p0_outen [1]),
    .opad(P0[1]));  // ../RTL/cmsdk_mcu_pin_mux.v(127)
  // ../RTL/cortexm0ds_logic.v(18793)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1092|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoax6_reg  (
    .a({_al_u1088_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .b({_al_u1089_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({_al_u1090_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1091_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] }),
    .mi({open_n1311,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ,_al_u1090_o}),
    .q({open_n1327,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[4] }));  // ../RTL/cortexm0ds_logic.v(18793)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1093|_al_u5995  (
    .a({open_n1328,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 }),
    .b({open_n1329,_al_u607_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ,_al_u932_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [4],_al_u5995_o}));
  // ../RTL/cortexm0ds_logic.v(18844)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1098|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6rax6_reg  (
    .a({_al_u1094_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({_al_u1095_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1096_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1097_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] }),
    .mi({open_n1357,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 ,_al_u1094_o}),
    .q({open_n1373,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] }));  // ../RTL/cortexm0ds_logic.v(18844)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u110 (
    .do({open_n1375,open_n1376,open_n1377,\u_cmsdk_mcu/p0_out [0]}),
    .ts(\u_cmsdk_mcu/p0_outen [0]),
    .opad(P0[0]));  // ../RTL/cmsdk_mcu_pin_mux.v(126)
  // ../RTL/cortexm0ds_logic.v(18799)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1101|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipoax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] }),
    .mi({open_n1393,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1101_o,_al_u874_o}),
    .q({open_n1409,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[5] }));  // ../RTL/cortexm0ds_logic.v(18799)
  // ../RTL/cortexm0ds_logic.v(18827)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1104|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8qax6_reg  (
    .a({_al_u1100_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({_al_u1101_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1102_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1103_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] }),
    .mi({open_n1420,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ,_al_u1102_o}),
    .q({open_n1425,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] }));  // ../RTL/cortexm0ds_logic.v(18827)
  // ../RTL/cortexm0ds_logic.v(18946)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1108|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltwax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] }),
    .mi({open_n1436,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y41pw6 ,_al_u726_o}),
    .q({open_n1441,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[13] }));  // ../RTL/cortexm0ds_logic.v(18946)
  EG_PHY_PAD #(
    //.LOCATION("A8"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u111 (
    .ipad(SWCLKTCK),
    .di(SWCLKTCK_pad));  // ../RTL/M0demo.v(15)
  // ../RTL/cortexm0ds_logic.v(18843)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1110|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4rax6_reg  (
    .a({_al_u1106_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .b({_al_u1107_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y41pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] }),
    .mi({open_n1469,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 ,_al_u1106_o}),
    .q({open_n1474,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] }));  // ../RTL/cortexm0ds_logic.v(18843)
  // ../RTL/cortexm0ds_logic.v(18800)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1114|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hroax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] }),
    .mi({open_n1485,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1114_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha4pw6 }),
    .q({open_n1490,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[6] }));  // ../RTL/cortexm0ds_logic.v(18800)
  // ../RTL/cortexm0ds_logic.v(18931)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1115|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozvax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] }),
    .mi({open_n1501,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1115_o,_al_u839_o}),
    .q({open_n1506,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] }));  // ../RTL/cortexm0ds_logic.v(18931)
  // ../RTL/cortexm0ds_logic.v(18828)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1116|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaqax6_reg  (
    .a({_al_u1112_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({_al_u1113_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1114_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1115_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] }),
    .mi({open_n1517,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ,_al_u1112_o}),
    .q({open_n1522,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[6] }));  // ../RTL/cortexm0ds_logic.v(18828)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u112 (
    .ipad(TDI));  // ../RTL/M0demo.v(12)
  // ../RTL/cortexm0ds_logic.v(18945)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1120|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrwax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] }),
    .mi({open_n1551,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0pw6 ,_al_u731_o}),
    .q({open_n1556,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[14] }));  // ../RTL/cortexm0ds_logic.v(18945)
  // ../RTL/cortexm0ds_logic.v(18917)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1122|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V7vax6_reg  (
    .a({_al_u1118_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({_al_u1119_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1121_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] }),
    .mi({open_n1560,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 ,_al_u1119_o}),
    .q({open_n1576,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] }));  // ../RTL/cortexm0ds_logic.v(18917)
  // ../RTL/cortexm0ds_logic.v(18932)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1125|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N1wax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] }),
    .mi({open_n1587,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u1125_o,_al_u888_o}),
    .q({open_n1592,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[7] }));  // ../RTL/cortexm0ds_logic.v(18932)
  // ../RTL/cortexm0ds_logic.v(18829)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1128|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wcqax6_reg  (
    .a({_al_u1124_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({_al_u1125_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1126_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc0pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] }),
    .mi({open_n1596,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ,_al_u1126_o}),
    .q({open_n1612,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] }));  // ../RTL/cortexm0ds_logic.v(18829)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u113 (
    .do({open_n1614,open_n1615,open_n1616,1'b0}),
    .ts(1'b1),
    .opad(TDO));  // ../RTL/cmsdk_mcu_pin_mux.v(211)
  // ../RTL/cortexm0ds_logic.v(19786)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1131|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zv7bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] }),
    .mi({open_n1632,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1131_o,_al_u737_o}),
    .q({open_n1648,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[15] }));  // ../RTL/cortexm0ds_logic.v(19786)
  // ../RTL/cortexm0ds_logic.v(19785)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1134|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt7bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .b({_al_u1131_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({_al_u1132_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1133_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] }),
    .mi({open_n1659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 ,_al_u1133_o}),
    .q({open_n1664,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] }));  // ../RTL/cortexm0ds_logic.v(19785)
  // ../RTL/cortexm0ds_logic.v(18943)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1136|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lnwax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] }),
    .mi({open_n1675,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzow6 ,_al_u750_o}),
    .q({open_n1680,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[17] }));  // ../RTL/cortexm0ds_logic.v(18943)
  EG_PHY_PAD #(
    //.LOCATION("K14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u114 (
    .ipad(XTAL1),
    .di(XTAL1_pad));  // ../RTL/M0demo.v(5)
  // ../RTL/cortexm0ds_logic.v(18840)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1140|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyqax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .b({_al_u1137_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1138_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1139_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] }),
    .mi({open_n1701,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 ,_al_u1139_o}),
    .q({open_n1717,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] }));  // ../RTL/cortexm0ds_logic.v(18840)
  // ../RTL/cortexm0ds_logic.v(18806)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1143|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3pax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] }),
    .mi({open_n1721,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({_al_u1143_o,_al_u766_o}),
    .q({open_n1737,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[1] }));  // ../RTL/cortexm0ds_logic.v(18806)
  // ../RTL/cortexm0ds_logic.v(18834)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1146|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmqax6_reg  (
    .a({_al_u1142_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({_al_u1143_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1144_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1145_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] }),
    .mi({open_n1748,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ,_al_u1144_o}),
    .q({open_n1753,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] }));  // ../RTL/cortexm0ds_logic.v(18834)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u1147|_al_u5989  (
    .a({open_n1754,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 }),
    .b({open_n1755,_al_u607_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ,_al_u932_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u115 (
    .do({open_n1777,open_n1778,open_n1779,XTAL2_pad}),
    .opad(XTAL2));  // ../RTL/M0demo.v(6)
  // ../RTL/cortexm0ds_logic.v(18801)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1150|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gtoax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] }),
    .mi({open_n1796,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u1150_o,_al_u1124_o}),
    .q({open_n1812,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] }));  // ../RTL/cortexm0ds_logic.v(18801)
  // ../RTL/cortexm0ds_logic.v(18839)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1152|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwqax6_reg  (
    .a({_al_u1148_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({_al_u1149_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1150_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] }),
    .mi({open_n1823,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 ,_al_u1149_o}),
    .q({open_n1828,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] }));  // ../RTL/cortexm0ds_logic.v(18839)
  // ../RTL/cortexm0ds_logic.v(18838)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1158|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uuqax6_reg  (
    .a({_al_u1154_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({_al_u1155_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1156_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1157_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] }),
    .mi({open_n1832,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 ,_al_u1157_o}),
    .q({open_n1848,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] }));  // ../RTL/cortexm0ds_logic.v(18838)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u116 (
    .do({open_n1850,open_n1851,open_n1852,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]),
    .di(b_pad_gpio_porta_pad[7]),
    .bpad(b_pad_gpio_porta[7]));  // ../RTL/gpio.v(182)
  // ../RTL/cortexm0ds_logic.v(18809)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1162|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9pax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] }),
    .mi({open_n1867,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .f({_al_u1162_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L27pw6 }),
    .q({open_n1883,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[20] }));  // ../RTL/cortexm0ds_logic.v(18809)
  // ../RTL/cortexm0ds_logic.v(18808)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1169|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E7pax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] }),
    .mi({open_n1887,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .f({_al_u1169_o,_al_u777_o}),
    .q({open_n1903,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[21] }));  // ../RTL/cortexm0ds_logic.v(18808)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u117 (
    .do({open_n1905,open_n1906,open_n1907,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]),
    .di(b_pad_gpio_porta_pad[6]),
    .bpad(b_pad_gpio_porta[6]));  // ../RTL/gpio.v(178)
  // ../RTL/cortexm0ds_logic.v(18836)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1170|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqqax6_reg  (
    .a({_al_u1166_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({_al_u1167_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1168_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1169_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] }),
    .mi({open_n1922,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 ,_al_u1167_o}),
    .q({open_n1938,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] }));  // ../RTL/cortexm0ds_logic.v(18836)
  // ../RTL/cortexm0ds_logic.v(19999)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1176|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Trebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({_al_u1173_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1174_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1175_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] }),
    .mi({open_n1942,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 ,_al_u1173_o}),
    .q({open_n1958,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] }));  // ../RTL/cortexm0ds_logic.v(19999)
  // ../RTL/cortexm0ds_logic.v(18822)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1179|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azpax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] }),
    .mi({open_n1969,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u1179_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Za6pw6 }),
    .q({open_n1974,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[23] }));  // ../RTL/cortexm0ds_logic.v(18822)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u118 (
    .do({open_n1976,open_n1977,open_n1978,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]),
    .di(b_pad_gpio_porta_pad[5]),
    .bpad(b_pad_gpio_porta[5]));  // ../RTL/gpio.v(174)
  // ../RTL/cortexm0ds_logic.v(18067)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1181|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv6ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] }),
    .mi({open_n2000,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u1181_o,_al_u792_o}),
    .q({open_n2005,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[23] }));  // ../RTL/cortexm0ds_logic.v(18067)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u1182|_al_u3604  (
    .a({_al_u1178_o,open_n2006}),
    .b({_al_u1179_o,open_n2007}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yow6 ,_al_u3603_o}),
    .d({_al_u1181_o,_al_u3601_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 }));
  // ../RTL/cortexm0ds_logic.v(18830)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1188|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veqax6_reg  (
    .a({_al_u1184_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({_al_u1185_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1186_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1187_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] }),
    .mi({open_n2031,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 ,_al_u1185_o}),
    .q({open_n2047,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] }));  // ../RTL/cortexm0ds_logic.v(18830)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u119 (
    .do({open_n2049,open_n2050,open_n2051,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]),
    .di(b_pad_gpio_porta_pad[4]),
    .bpad(b_pad_gpio_porta[4]));  // ../RTL/gpio.v(170)
  // ../RTL/cortexm0ds_logic.v(17933)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1192|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P21qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] }),
    .mi({open_n2066,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlxow6 ,_al_u879_o}),
    .q({open_n2082,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] }));  // ../RTL/cortexm0ds_logic.v(17933)
  // ../RTL/cortexm0ds_logic.v(18847)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1194|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcrax6_reg  (
    .a({_al_u1190_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkxow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlxow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1193_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] }),
    .mi({open_n2093,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkxow6 }),
    .q({open_n2098,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] }));  // ../RTL/cortexm0ds_logic.v(18847)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u120 (
    .do({open_n2100,open_n2101,open_n2102,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]),
    .di(b_pad_gpio_porta_pad[3]),
    .bpad(b_pad_gpio_porta[3]));  // ../RTL/gpio.v(166)
  // ../RTL/cortexm0ds_logic.v(18835)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1200|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoqax6_reg  (
    .a({_al_u1196_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .b({_al_u1197_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1198_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oaxow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] }),
    .mi({open_n2124,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oaxow6 }),
    .q({open_n2129,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] }));  // ../RTL/cortexm0ds_logic.v(18835)
  // ../RTL/cortexm0ds_logic.v(18818)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1202|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erpax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] }),
    .mi({open_n2140,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({_al_u1202_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D14pw6 }),
    .q({open_n2145,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[9] }));  // ../RTL/cortexm0ds_logic.v(18818)
  // ../RTL/cortexm0ds_logic.v(17946)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1203|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir1qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] }),
    .mi({open_n2156,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({_al_u1203_o,_al_u843_o}),
    .q({open_n2161,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[9] }));  // ../RTL/cortexm0ds_logic.v(17946)
  // ../RTL/cortexm0ds_logic.v(18846)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1206|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uarax6_reg  (
    .a({_al_u1202_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({_al_u1203_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1204_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] }),
    .mi({open_n2172,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 ,_al_u1204_o}),
    .q({open_n2177,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[9] }));  // ../RTL/cortexm0ds_logic.v(18846)
  // ../RTL/cortexm0ds_logic.v(18803)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1209|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fxoax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] }),
    .mi({open_n2188,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u1209_o,_al_u808_o}),
    .q({open_n2193,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[26] }));  // ../RTL/cortexm0ds_logic.v(18803)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u121 (
    .do({open_n2195,open_n2196,open_n2197,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]),
    .di(b_pad_gpio_porta_pad[2]),
    .bpad(b_pad_gpio_porta[2]));  // ../RTL/gpio.v(162)
  // ../RTL/cortexm0ds_logic.v(17692)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1212|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvtpw6_reg  (
    .a({_al_u1208_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .b({_al_u1209_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1210_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1211_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] }),
    .mi({open_n2219,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 ,_al_u1210_o}),
    .q({open_n2224,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[26] }));  // ../RTL/cortexm0ds_logic.v(17692)
  // ../RTL/cortexm0ds_logic.v(17537)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1216|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfppw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] }),
    .mi({open_n2228,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u1216_o,_al_u814_o}),
    .q({open_n2244,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[27] }));  // ../RTL/cortexm0ds_logic.v(17537)
  // ../RTL/cortexm0ds_logic.v(18907)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1218|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnuax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjwow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({_al_u1215_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({_al_u1216_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1217_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] }),
    .mi({open_n2248,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 ,_al_u1215_o}),
    .q({open_n2264,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] }));  // ../RTL/cortexm0ds_logic.v(18907)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u122 (
    .do({open_n2266,open_n2267,open_n2268,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [1]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]),
    .di(b_pad_gpio_porta_pad[1]),
    .bpad(b_pad_gpio_porta[1]));  // ../RTL/gpio.v(158)
  // ../RTL/cortexm0ds_logic.v(20175)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1222|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] }),
    .mi({open_n2283,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9wow6 ,_al_u821_o}),
    .q({open_n2299,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[28] }));  // ../RTL/cortexm0ds_logic.v(20175)
  // ../RTL/cortexm0ds_logic.v(20168)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1223|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9ibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] }),
    .mi({open_n2310,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({_al_u1223_o,_al_u822_o}),
    .q({open_n2315,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[28] }));  // ../RTL/cortexm0ds_logic.v(20168)
  // ../RTL/cortexm0ds_logic.v(20174)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1224|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlibx6_reg  (
    .a({_al_u1220_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .b({_al_u1221_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9wow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1223_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] }),
    .mi({open_n2319,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 ,_al_u1220_o}),
    .q({open_n2335,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] }));  // ../RTL/cortexm0ds_logic.v(20174)
  // ../RTL/cortexm0ds_logic.v(18926)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1229|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rpvax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] }),
    .mi({open_n2339,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({_al_u1229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4pw6 }),
    .q({open_n2355,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[30] }));  // ../RTL/cortexm0ds_logic.v(18926)
  EG_PHY_PAD #(
    //.LOCATION("N3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .TSMUX("INV"))
    _al_u123 (
    .do({open_n2357,open_n2358,open_n2359,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [0]}),
    .ts(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]),
    .di(b_pad_gpio_porta_pad[0]),
    .bpad(b_pad_gpio_porta[0]));  // ../RTL/gpio.v(154)
  // ../RTL/cortexm0ds_logic.v(17201)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1230|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Weipw6_reg  (
    .a({_al_u1226_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({_al_u1227_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({_al_u1228_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] }),
    .mi({open_n2374,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 ,_al_u1226_o}),
    .q({open_n2390,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] }));  // ../RTL/cortexm0ds_logic.v(17201)
  // ../RTL/cortexm0ds_logic.v(18796)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1236|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjoax6_reg  (
    .a({_al_u1232_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .b({_al_u1233_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({_al_u1234_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1235_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] }),
    .mi({open_n2401,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 ,_al_u1233_o}),
    .q({open_n2406,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] }));  // ../RTL/cortexm0ds_logic.v(18796)
  // ../RTL/cortexm0ds_logic.v(19721)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1238|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No5bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] }),
    .mi({open_n2417,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u1238_o,_al_u828_o}),
    .q({open_n2422,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[29] }));  // ../RTL/cortexm0ds_logic.v(19721)
  EG_PHY_PAD #(
    //.LOCATION("R5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u124 (
    .ipad(nTRST));  // ../RTL/M0demo.v(11)
  // ../RTL/cortexm0ds_logic.v(18805)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1240|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1pax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] }),
    .mi({open_n2451,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u1240_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4pw6 }),
    .q({open_n2456,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[29] }));  // ../RTL/cortexm0ds_logic.v(18805)
  // ../RTL/cortexm0ds_logic.v(18936)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1242|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M9wax6_reg  (
    .a({_al_u1238_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({_al_u1239_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1240_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1241_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] }),
    .mi({open_n2467,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 ,_al_u1239_o}),
    .q({open_n2472,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] }));  // ../RTL/cortexm0ds_logic.v(18936)
  // ../RTL/cortexm0ds_logic.v(18813)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1246|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehpax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] }),
    .mi({open_n2476,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .f({_al_u1246_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad8pw6 }),
    .q({open_n2492,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[16] }));  // ../RTL/cortexm0ds_logic.v(18813)
  // ../RTL/cortexm0ds_logic.v(18944)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1248|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lpwax6_reg  (
    .a({_al_u1244_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({_al_u1245_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({_al_u1246_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1247_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] }),
    .mi({open_n2496,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 ,_al_u1245_o}),
    .q({open_n2512,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] }));  // ../RTL/cortexm0ds_logic.v(18944)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u125 (
    .do({open_n2514,open_n2515,open_n2516,uart0_txd_pad}),
    .opad(uart0_txd));  // ../RTL/M0demo.v(20)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1251|_al_u3256  (
    .b({open_n2532,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .f({_al_u1251_o,_al_u3256_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1252|_al_u1250  (
    .b({_al_u1251_o,open_n2559}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({_al_u1250_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ,_al_u1250_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1255|_al_u1256  (
    .b({open_n2582,_al_u1255_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ,_al_u1253_o}),
    .f({_al_u1255_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U73iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1257|_al_u903  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u903_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u1257_o,_al_u903_o}));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u126 (
    .do({open_n2636,open_n2637,open_n2638,uart0_txen_pad}),
    .opad(uart0_txen));  // ../RTL/M0demo.v(21)
  // ../RTL/cmsdk_apb_uart.v(392)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1260|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u467_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n50 ),
    .clk(XTAL1_wire),
    .d({_al_u473_o,_al_u473_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 }),
    .q({open_n2673,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full }));  // ../RTL/cmsdk_apb_uart.v(392)
  // ../RTL/cmsdk_apb_uart.v(220)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D*~(C*A)))"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("~(~B*~(D*~(C*A)))"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111111001100),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1101111111001100),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1261|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun_reg  (
    .a({open_n2674,\u_cmsdk_mcu/HWDATA [3]}),
    .b({open_n2675,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n17 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n17 ,open_n2692}),
    .q({open_n2696,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun }));  // ../RTL/cmsdk_apb_uart.v(220)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1263|_al_u681  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,_al_u681_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~(D*B*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000011100001111),
    .MODE("LOGIC"))
    \_al_u1265|_al_u606  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,open_n2721}),
    .b({_al_u606_o,open_n2722}),
    .c({_al_u1264_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 ,_al_u606_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1267|_al_u1266  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ,_al_u1266_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1269|_al_u2862  (
    .b({open_n2773,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,_al_u2861_o}),
    .f({_al_u1269_o,_al_u2862_o}));
  // ../RTL/cortexm0ds_logic.v(18730)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~C*~B*A)"),
    //.LUTF1("(A*~(~C*~(D*B)))"),
    //.LUTG0("~(D*~C*~B*A)"),
    //.LUTG1("(A*~(~C*~(D*B)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110111111111),
    .INIT_LUTF1(16'b1010100010100000),
    .INIT_LUTG0(16'b1111110111111111),
    .INIT_LUTG1(16'b1010100010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1270|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6_reg  (
    .a({_al_u1268_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 }),
    .b({_al_u1269_o,_al_u1270_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,_al_u1273_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1270_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 }),
    .q({open_n2817,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 }));  // ../RTL/cortexm0ds_logic.v(18730)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1272|_al_u1271  (
    .c({_al_u1271_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u1269_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ,_al_u1271_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*B*~(~D*~A))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1100000010000000),
    .MODE("LOGIC"))
    \_al_u1273|_al_u604  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ,open_n2842}),
    .b({_al_u604_o,open_n2843}),
    .c({_al_u609_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u1273_o,_al_u604_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1275|_al_u1274  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~B*~(~D*C*A))"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~B*~(~D*C*A))"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0011001100010011),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0011001100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1277|_al_u1276  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ,_al_u681_o}),
    .b({_al_u1276_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u682_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 ,_al_u1276_o}));
  // ../RTL/cmsdk_apb_uart.v(229)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D*~(C*A)))"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("~(~B*~(D*~(C*A)))"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111111001100),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1101111111001100),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1280|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun_reg  (
    .a({open_n2912,\u_cmsdk_mcu/HWDATA [2]}),
    .b({open_n2913,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n9_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n20 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n20 ,open_n2930}),
    .q({open_n2934,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun }));  // ../RTL/cmsdk_apb_uart.v(229)
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1281|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b7  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [8],_al_u4237_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u1281_o,\u_cmsdk_mcu/HADDR [9]}),
    .q({open_n2957,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [7]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1282|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8],open_n2958}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4],_al_u4141_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u1282_o,\u_cmsdk_mcu/HADDR [6]}),
    .q({open_n2975,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1283|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b2  (
    .a({_al_u1281_o,open_n2976}),
    .b({_al_u1282_o,_al_u4231_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1],\u_cmsdk_mcu/HADDR [4]}),
    .q({open_n2997,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1284|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0],_al_u4225_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],\u_cmsdk_mcu/HADDR [3]}),
    .q({open_n3016,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  // ../RTL/cortexm0ds_logic.v(19095)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1285|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6_reg  (
    .a({\u_cmsdk_mcu/sram_hrdata [30],open_n3017}),
    .b({\u_cmsdk_mcu/flash_hrdata [30],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/flash_hrdata [30]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/HWDATA [30]}),
    .mi({open_n3028,\u_cmsdk_mcu/HWDATA [30]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1285_o,\u_cmsdk_mcu/u_ahb_rom/n13 [30]}),
    .q({open_n3032,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 }));  // ../RTL/cortexm0ds_logic.v(19095)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1286|_al_u1865  (
    .c({_al_u1285_o,_al_u1864_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]}),
    .f({_al_u1286_o,_al_u1865_o}));
  // ../RTL/cortexm0ds_logic.v(17690)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1288|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ,open_n3061}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [10]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ,_al_u2339_o}),
    .f({_al_u1288_o,open_n3076}),
    .q({open_n3080,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 }));  // ../RTL/cortexm0ds_logic.v(17690)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1289|_al_u6675  (
    .a({_al_u1288_o,_al_u6673_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ,_al_u6674_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 }),
    .f({_al_u1289_o,_al_u6675_o}));
  // ../RTL/cortexm0ds_logic.v(17928)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1290|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ,open_n3105}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [8]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ,_al_u2343_o}),
    .f({_al_u1290_o,open_n3124}),
    .q({open_n3128,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 }));  // ../RTL/cortexm0ds_logic.v(17928)
  // ../RTL/cortexm0ds_logic.v(18962)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1291|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ,open_n3129}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [14]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ,_al_u2331_o}),
    .f({_al_u1291_o,open_n3148}),
    .q({open_n3152,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 }));  // ../RTL/cortexm0ds_logic.v(18962)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1292|_al_u1294  (
    .a({open_n3153,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 }),
    .b({_al_u1290_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 }),
    .c({_al_u1291_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 }),
    .d({_al_u1289_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 }),
    .f({_al_u1292_o,_al_u1294_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1293|_al_u5367  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ,_al_u5067_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 }),
    .f({_al_u1293_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dooow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1295|_al_u5984  (
    .b({_al_u1293_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 }),
    .c({_al_u1294_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] }),
    .d({_al_u1292_o,_al_u5983_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ,_al_u5984_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u1296|_al_u2387  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u1296_o,_al_u2387_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1297|_al_u905  (
    .b({_al_u1296_o,open_n3250}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u1297_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u1299|_al_u1298  (
    .b({_al_u604_o,open_n3273}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u1297_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u1299_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*~A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000010000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1300|_al_u4488  (
    .a({open_n3294,_al_u4485_o}),
    .b({open_n3295,_al_u1299_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 ,_al_u1777_o}),
    .d({_al_u1299_o,_al_u4487_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ,_al_u4488_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1301|_al_u2311  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 }),
    .f({_al_u1301_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1302|_al_u578  (
    .b({open_n3340,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(20225)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*~(~D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100110001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1305|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ,open_n3365}),
    .b({_al_u1304_o,open_n3366}),
    .c({_al_u405_o,_al_u1305_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,_al_u1301_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1305_o,open_n3380}),
    .q({open_n3384,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 }));  // ../RTL/cortexm0ds_logic.v(20225)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(C@(D*A)))"),
    //.LUT1("(~B*(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT_LUT0(16'b0001001000110000),
    .INIT_LUT1(16'b0011000000010001),
    .MODE("LOGIC"))
    \_al_u1307|_al_u530  (
    .a({_al_u530_o,_al_u529_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .f({_al_u1307_o,_al_u530_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*~D))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~B*~(~C*~D))"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0011001100110000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0011001100110000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1310|_al_u1309  (
    .b({_al_u1309_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .d({_al_u1250_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .f({_al_u1310_o,_al_u1309_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1311|_al_u1308  (
    .a({_al_u1308_o,open_n3431}),
    .b({_al_u1310_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .c({_al_u1251_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ,_al_u1250_o}),
    .f({_al_u1311_o,_al_u1308_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(A*~(~D*~(~C*B)))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(A*~(~D*~(~C*B)))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1010101000001000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1010101000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1313|_al_u1312  (
    .a({_al_u1307_o,open_n3456}),
    .b({_al_u1311_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ,_al_u529_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tw2iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(D*~C*B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"))
    \_al_u1315|_al_u713  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(18771)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1316|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S5nax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] }),
    .mi({open_n3504,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({_al_u1316_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qy2pw6 }),
    .q({open_n3520,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[0] }));  // ../RTL/cortexm0ds_logic.v(18771)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*~A)"),
    //.LUT1("(~D*~C*B*A)"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"))
    \_al_u1317|_al_u710  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*A)"),
    //.LUTF1("(~D*~C*B*~A)"),
    //.LUTG0("(D*~C*~B*A)"),
    //.LUTG1("(~D*~C*B*~A)"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1318|_al_u707  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~A)"),
    //.LUTF1("(D*C*B*~A)"),
    //.LUTG0("(D*~C*~B*~A)"),
    //.LUTG1("(D*C*B*~A)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b0000000100000000),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1320|_al_u706  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(18853)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1323|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qorax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .b({_al_u1316_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .c({_al_u1319_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls9pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] }),
    .mi({open_n3599,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({_al_u1323_o,_al_u1319_o}),
    .q({open_n3604,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] }));  // ../RTL/cortexm0ds_logic.v(18853)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1326|_al_u1325  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u1327|_al_u914  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ,open_n3633}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ,open_n3634}),
    .c({_al_u914_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u1271_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u1327_o,_al_u914_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*~A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000010000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u1328|_al_u1321  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 }),
    .f({_al_u1328_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~D*~(C*~B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1331|_al_u1330  (
    .b({_al_u1329_o,open_n3677}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u1328_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u1331_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1334|_al_u1333  (
    .a({_al_u1327_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .b({_al_u1331_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u1332_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u1333_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u1334_o,_al_u1333_o}));
  // ../RTL/cortexm0ds_logic.v(17324)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*A*~(D*B))"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("~(~C*A*~(D*B))"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110111110101),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b1111110111110101),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1335|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6_reg  (
    .a({open_n3726,_al_u4212_o}),
    .b({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ,_al_u4213_o}),
    .clk(XTAL1_wire),
    .d({_al_u1323_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ,open_n3745}),
    .q({open_n3749,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 }));  // ../RTL/cortexm0ds_logic.v(17324)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u1337|_al_u1336  (
    .b({_al_u1336_o,open_n3752}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u1337_o,_al_u1336_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1339|_al_u1338  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ,open_n3775}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u1337_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u1339_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~B*A)"),
    //.LUTF1("(~A*~(~D*~(~C*~B)))"),
    //.LUTG0("(D*C*~B*A)"),
    //.LUTG1("(~A*~(~D*~(~C*~B)))"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0101010100000001),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0101010100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1343|_al_u1341  (
    .a({_al_u1341_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u1342_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u1343_o,_al_u1341_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("~(A*~((C*B))*~(D)+A*(C*B)*~(D)+~(A)*(C*B)*D+A*(C*B)*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("~(A*~((C*B))*~(D)+A*(C*B)*~(D)+~(A)*(C*B)*D+A*(C*B)*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0011111101010101),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0011111101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1345|_al_u696  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ,open_n3824}),
    .b({_al_u696_o,open_n3825}),
    .c({_al_u1344_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u1345_o,_al_u696_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~A*~(~D*C)))"),
    //.LUT1("(~D*C*B*A)"),
    .INIT_LUT0(16'b0010001000110010),
    .INIT_LUT1(16'b0000000010000000),
    .MODE("LOGIC"))
    \_al_u1348|_al_u1347  (
    .a({_al_u1339_o,_al_u1346_o}),
    .b({_al_u1343_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({_al_u1345_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u1347_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u1348_o,_al_u1347_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1349|_al_u1617  (
    .c({_al_u1348_o,_al_u1348_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ,_al_u1616_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [7]}));
  // ../RTL/cortexm0ds_logic.v(20171)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1351|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] }),
    .mi({open_n3908,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({_al_u1351_o,_al_u1519_o}),
    .q({open_n3913,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] }));  // ../RTL/cortexm0ds_logic.v(20171)
  // ../RTL/cortexm0ds_logic.v(17884)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1352|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Onypw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] }),
    .mi({open_n3917,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87pw6 ,_al_u1967_o}),
    .q({open_n3933,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[1] }));  // ../RTL/cortexm0ds_logic.v(17884)
  // ../RTL/cortexm0ds_logic.v(17882)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1353|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjypw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1350_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1351_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] }),
    .mi({open_n3937,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V77pw6 ,_al_u1350_o}),
    .q({open_n3953,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[1] }));  // ../RTL/cortexm0ds_logic.v(17882)
  // ../RTL/cortexm0ds_logic.v(18854)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1354|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqrax6_reg  (
    .a({open_n3954,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V77pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] }),
    .mi({open_n3958,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({_al_u1354_o,_al_u1964_o}),
    .q({open_n3974,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[1] }));  // ../RTL/cortexm0ds_logic.v(18854)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1355|_al_u1609  (
    .c({_al_u1348_o,_al_u1348_o}),
    .d({_al_u1354_o,_al_u1608_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [8]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1358|_al_u1357  (
    .a({open_n4003,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .b({open_n4004,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({_al_u1357_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ,_al_u1357_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u1360|_al_u1359  (
    .b({_al_u1359_o,open_n4027}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u1360_o,_al_u1359_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1362|_al_u3682  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1363|_al_u1799  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv }),
    .f({_al_u1363_o,_al_u1799_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(~D*C)))"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1000100011001000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u1364|_al_u4158  (
    .a({open_n4100,_al_u4157_o}),
    .b({_al_u1363_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({_al_u1364_o,_al_u4158_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(~(B)*C*~(D)+B*~(C)*D+B*C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b1000100000100000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u1365|_al_u1361  (
    .a({open_n4121,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv }),
    .b({_al_u1364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B91ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 }));
  // ../RTL/cortexm0ds_logic.v(17279)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(B*~(C*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1366|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6_reg  (
    .a({open_n4142,_al_u1366_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B91ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ),
    .clk(XTAL1_wire),
    .d({_al_u1360_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 }),
    .f({_al_u1366_o,open_n4160}),
    .q({open_n4164,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 }));  // ../RTL/cortexm0ds_logic.v(17279)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1010111100110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1010111100110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1372|_al_u1649  (
    .a({open_n4165,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u1359_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u1372_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8aiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(~D*~B*~(~C*A))"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(~D*~B*~(~C*A))"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b0000000000110001),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000000000110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1373|_al_u1368  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ,open_n4190}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ,_al_u1367_o}),
    .c({_al_u1370_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u1372_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~(A)*C*~(D)+A*C*~(D)+~(A)*~(C)*D+A*~(C)*D+A*C*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*(~(A)*C*~(D)+A*C*~(D)+~(A)*~(C)*D+A*~(C)*D+A*C*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0010001100110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0010001100110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1374|_al_u3681  (
    .a({open_n4215,_al_u3679_o}),
    .b({open_n4216,_al_u3680_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ,_al_u3681_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000100110001),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0000000100110001),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1377|_al_u1376  (
    .a({open_n4241,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .b({_al_u1375_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({_al_u1376_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ,_al_u1376_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B*~(C*A)))"),
    //.LUTF1("(~B*A*~(D*C))"),
    //.LUTG0("(D*~(B*~(C*A)))"),
    //.LUTG1("(~B*A*~(D*C))"),
    .INIT_LUTF0(16'b1011001100000000),
    .INIT_LUTF1(16'b0000001000100010),
    .INIT_LUTG0(16'b1011001100000000),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1379|_al_u917  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .b({_al_u908_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u1379_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1380|_al_u3214  (
    .a({_al_u912_o,open_n4290}),
    .b({_al_u696_o,open_n4291}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({_al_u1380_o,_al_u3214_o}));
  // ../RTL/cortexm0ds_logic.v(17848)
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("~(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110111010101),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1101110111010101),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1381|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6_reg  (
    .a({_al_u1379_o,_al_u1381_o}),
    .b({_al_u1380_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ,_al_u1382_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ,_al_u1383_o}),
    .f({_al_u1381_o,open_n4333}),
    .q({open_n4337,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }));  // ../RTL/cortexm0ds_logic.v(17848)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u1382|_al_u3602  (
    .a({open_n4338,_al_u3120_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 }),
    .d({_al_u916_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 }),
    .f({_al_u1382_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqniu6 }));
  // ../RTL/cortexm0ds_logic.v(18337)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*C)*~(B*A))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("~(~(D*C)*~(B*A))"),
    //.LUTG1("(D*C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111100010001000),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b1111100010001000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1387|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u1387_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u1387_o,open_n4376}),
    .q({open_n4380,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 }));  // ../RTL/cortexm0ds_logic.v(18337)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1389|_al_u1392  (
    .a({_al_u702_o,_al_u702_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 }));
  // ../RTL/cortexm0ds_logic.v(17924)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1390|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tk0qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,open_n4405}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,_al_u1390_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 }),
    .mi({open_n4409,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u1390_o,_al_u1391_o}),
    .q({open_n4425,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] }));  // ../RTL/cortexm0ds_logic.v(17924)
  // ../RTL/cortexm0ds_logic.v(17233)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1393|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bdjpw6_reg  (
    .a({open_n4426,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1391_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[10] }),
    .mi({open_n4437,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u1393_o,_al_u2081_o}),
    .q({open_n4442,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[10] }));  // ../RTL/cortexm0ds_logic.v(17233)
  // ../RTL/cortexm0ds_logic.v(18892)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1395|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eutax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] }),
    .mi({open_n4446,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u1395_o,_al_u2080_o}),
    .q({open_n4462,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[12] }));  // ../RTL/cortexm0ds_logic.v(18892)
  // ../RTL/cortexm0ds_logic.v(18789)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1396|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5oax6_reg  (
    .a({open_n4463,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1394_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .c({_al_u1395_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1393_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] }),
    .mi({open_n4474,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u1396_o,_al_u1394_o}),
    .q({open_n4479,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[12] }));  // ../RTL/cortexm0ds_logic.v(18789)
  // ../RTL/cortexm0ds_logic.v(17531)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1397|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O3ppw6_reg  (
    .a({_al_u1396_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] }),
    .mi({open_n4490,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u1397_o,_al_u2078_o}),
    .q({open_n4495,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[12] }));  // ../RTL/cortexm0ds_logic.v(17531)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100010011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1398|_al_u5932  (
    .a({open_n4496,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 }),
    .b({open_n4497,_al_u5931_o}),
    .c({_al_u1348_o,_al_u1397_o}),
    .d({_al_u1397_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [12],_al_u5932_o}));
  // ../RTL/cortexm0ds_logic.v(18863)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1399|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8sax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] }),
    .mi({open_n4528,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({_al_u1399_o,_al_u2104_o}),
    .q({open_n4533,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[13] }));  // ../RTL/cortexm0ds_logic.v(18863)
  // ../RTL/cortexm0ds_logic.v(17923)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1400|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ti0qw6_reg  (
    .a({open_n4534,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({_al_u1399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] }),
    .mi({open_n4538,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({_al_u1400_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0pw6 }),
    .q({open_n4554,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[11] }));  // ../RTL/cortexm0ds_logic.v(17923)
  // ../RTL/cortexm0ds_logic.v(18788)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1403|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3oax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 }),
    .mi({open_n4565,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({_al_u1403_o,_al_u2102_o}),
    .q({open_n4570,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[13] }));  // ../RTL/cortexm0ds_logic.v(18788)
  // ../RTL/cortexm0ds_logic.v(17302)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1404|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnkpw6_reg  (
    .b({_al_u1402_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 }),
    .c({_al_u1403_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1401_o,_al_u1400_o}),
    .mi({open_n4583,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({_al_u1404_o,_al_u1401_o}),
    .q({open_n4588,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[11] }));  // ../RTL/cortexm0ds_logic.v(17302)
  // ../RTL/cortexm0ds_logic.v(18967)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1405|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6_reg  (
    .a({_al_u1404_o,open_n4589}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ,_al_u4128_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 ,_al_u4126_o}),
    .f({_al_u1405_o,open_n4604}),
    .q({open_n4608,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 }));  // ../RTL/cortexm0ds_logic.v(18967)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100010011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1406|_al_u5953  (
    .a({open_n4609,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 }),
    .b({open_n4610,_al_u5952_o}),
    .c({_al_u1348_o,_al_u1405_o}),
    .d({_al_u1405_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [13],_al_u5953_o}));
  // ../RTL/cortexm0ds_logic.v(18760)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1407|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjmax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,open_n4631}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,_al_u7010_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] ,_al_u6193_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] ,_al_u6969_o}),
    .f({_al_u1407_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .q({open_n4648,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] }));  // ../RTL/cortexm0ds_logic.v(18760)
  // ../RTL/cortexm0ds_logic.v(18117)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1408|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S78ax6_reg  (
    .a({open_n4649,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({_al_u1407_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] }),
    .mi({open_n4660,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({_al_u1408_o,_al_u2126_o}),
    .q({open_n4665,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[12] }));  // ../RTL/cortexm0ds_logic.v(18117)
  // ../RTL/cortexm0ds_logic.v(18114)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1410|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[14] }),
    .mi({open_n4676,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({_al_u1410_o,_al_u2122_o}),
    .q({open_n4681,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[14] }));  // ../RTL/cortexm0ds_logic.v(18114)
  // ../RTL/cortexm0ds_logic.v(18862)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1411|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O6sax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 }),
    .mi({open_n4692,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({_al_u1411_o,_al_u2124_o}),
    .q({open_n4697,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[14] }));  // ../RTL/cortexm0ds_logic.v(18862)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1412|_al_u6870  (
    .b({_al_u1410_o,open_n4700}),
    .c({_al_u1411_o,_al_u6869_o}),
    .d({_al_u1409_o,_al_u6868_o}),
    .f({_al_u1412_o,_al_u6870_o}));
  // ../RTL/cortexm0ds_logic.v(18119)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1413|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6_reg  (
    .a({_al_u1412_o,open_n4721}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ,_al_u4133_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ,_al_u4131_o}),
    .f({_al_u1413_o,open_n4740}),
    .q({open_n4744,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 }));  // ../RTL/cortexm0ds_logic.v(18119)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*B*~A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1011000011110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1414|_al_u6192  (
    .a({open_n4745,_al_u1413_o}),
    .b({open_n4746,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 }),
    .c({_al_u1348_o,_al_u6191_o}),
    .d({_al_u1413_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [14],_al_u6192_o}));
  // ../RTL/cortexm0ds_logic.v(19790)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1415|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z38bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] }),
    .mi({open_n4770,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1415_o,_al_u2146_o}),
    .q({open_n4786,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[15] }));  // ../RTL/cortexm0ds_logic.v(19790)
  // ../RTL/cortexm0ds_logic.v(19798)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1417|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zj8bx6_reg  (
    .a({open_n4787,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1416_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] }),
    .mi({open_n4798,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1417_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00pw6 }),
    .q({open_n4803,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[13] }));  // ../RTL/cortexm0ds_logic.v(19798)
  // ../RTL/cortexm0ds_logic.v(19791)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1418|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z58bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] }),
    .mi({open_n4814,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1418_o,_al_u2148_o}),
    .q({open_n4819,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[15] }));  // ../RTL/cortexm0ds_logic.v(19791)
  // ../RTL/cortexm0ds_logic.v(19797)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1420|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zh8bx6_reg  (
    .a({open_n4820,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1418_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .c({_al_u1419_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1417_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] }),
    .mi({open_n4831,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1420_o,_al_u1419_o}),
    .q({open_n4836,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[15] }));  // ../RTL/cortexm0ds_logic.v(19797)
  // ../RTL/cortexm0ds_logic.v(19796)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1421|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8bx6_reg  (
    .a({_al_u1420_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] }),
    .mi({open_n4847,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1421_o,_al_u2144_o}),
    .q({open_n4852,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[15] }));  // ../RTL/cortexm0ds_logic.v(19796)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100010011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1422|_al_u6177  (
    .a({open_n4853,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 }),
    .b({open_n4854,_al_u6176_o}),
    .c({_al_u1348_o,_al_u1421_o}),
    .d({_al_u1421_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [15],_al_u6177_o}));
  // ../RTL/cortexm0ds_logic.v(18786)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1423|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nznax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] }),
    .mi({open_n4885,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .f({_al_u1423_o,_al_u2283_o}),
    .q({open_n4890,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[16] }));  // ../RTL/cortexm0ds_logic.v(18786)
  // ../RTL/cortexm0ds_logic.v(17813)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1425|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfwpw6_reg  (
    .a({open_n4891,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1424_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] }),
    .mi({open_n4895,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .f({_al_u1425_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peqow6 }),
    .q({open_n4911,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[14] }));  // ../RTL/cortexm0ds_logic.v(17813)
  // ../RTL/cortexm0ds_logic.v(17811)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1426|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbwpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] }),
    .mi({open_n4915,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .f({_al_u1426_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ciqow6 }),
    .q({open_n4931,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[16] }));  // ../RTL/cortexm0ds_logic.v(17811)
  // ../RTL/cortexm0ds_logic.v(18889)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1427|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eotax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] }),
    .mi({open_n4942,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .f({_al_u1427_o,_al_u2285_o}),
    .q({open_n4947,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[16] }));  // ../RTL/cortexm0ds_logic.v(18889)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1428|_al_u745  (
    .a({open_n4948,_al_u741_o}),
    .b({_al_u1426_o,_al_u742_o}),
    .c({_al_u1427_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad8pw6 }),
    .d({_al_u1425_o,_al_u744_o}),
    .f({_al_u1428_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1429|_al_u746  (
    .a({_al_u1428_o,open_n4969}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ,open_n4970}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1429_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(D*~C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100010011001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100010011001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1430|_al_u5922  (
    .a({open_n4995,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 }),
    .b({open_n4996,_al_u5921_o}),
    .c({_al_u1348_o,_al_u1429_o}),
    .d({_al_u1429_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [16],_al_u5922_o}));
  // ../RTL/cortexm0ds_logic.v(17706)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1432|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydupw6_reg  (
    .a({open_n5021,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .b({_al_u1431_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] }),
    .mi({open_n5025,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u1432_o,_al_u1431_o}),
    .q({open_n5041,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] }));  // ../RTL/cortexm0ds_logic.v(17706)
  // ../RTL/cortexm0ds_logic.v(17921)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1433|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Te0qw6_reg  (
    .a({open_n5042,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1432_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] }),
    .mi({open_n5053,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u1433_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drzow6 }),
    .q({open_n5058,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[15] }));  // ../RTL/cortexm0ds_logic.v(17921)
  // ../RTL/cortexm0ds_logic.v(18785)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1435|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxnax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] }),
    .mi({open_n5062,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u1435_o,_al_u2165_o}),
    .q({open_n5078,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[17] }));  // ../RTL/cortexm0ds_logic.v(18785)
  // ../RTL/cortexm0ds_logic.v(17705)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1436|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ybupw6_reg  (
    .a({open_n5079,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({_al_u1435_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1433_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] }),
    .mi({open_n5090,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u1436_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18pw6 }),
    .q({open_n5095,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[17] }));  // ../RTL/cortexm0ds_logic.v(17705)
  // ../RTL/cortexm0ds_logic.v(19929)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1437|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6_reg  (
    .a({_al_u1436_o,open_n5096}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ,_al_u4063_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 ,_al_u4061_o}),
    .f({_al_u1437_o,open_n5111}),
    .q({open_n5115,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 }));  // ../RTL/cortexm0ds_logic.v(19929)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(D*~C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100010011001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100010011001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1438|_al_u6203  (
    .a({open_n5116,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 }),
    .b({open_n5117,_al_u6202_o}),
    .c({_al_u1348_o,_al_u1437_o}),
    .d({_al_u1437_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [17],_al_u6203_o}));
  // ../RTL/cortexm0ds_logic.v(18859)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1439|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O0sax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 }),
    .mi({open_n5145,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u1439_o,_al_u2204_o}),
    .q({open_n5161,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[18] }));  // ../RTL/cortexm0ds_logic.v(18859)
  // ../RTL/cortexm0ds_logic.v(17835)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1441|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pcxpw6_reg  (
    .a({open_n5162,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1440_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] }),
    .mi({open_n5173,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u1441_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eazow6 }),
    .q({open_n5178,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[16] }));  // ../RTL/cortexm0ds_logic.v(17835)
  // ../RTL/cortexm0ds_logic.v(18784)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1443|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvnax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] }),
    .mi({open_n5182,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u1443_o,_al_u2202_o}),
    .q({open_n5198,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[18] }));  // ../RTL/cortexm0ds_logic.v(18784)
  // ../RTL/cortexm0ds_logic.v(17832)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1444|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P6xpw6_reg  (
    .a({open_n5199,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs7pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({_al_u1443_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1441_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] }),
    .mi({open_n5203,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u1444_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs7pw6 }),
    .q({open_n5219,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[18] }));  // ../RTL/cortexm0ds_logic.v(17832)
  // ../RTL/cortexm0ds_logic.v(20214)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1445|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6_reg  (
    .a({_al_u1444_o,open_n5220}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ,_al_u4068_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 ,_al_u4066_o}),
    .f({_al_u1445_o,open_n5239}),
    .q({open_n5243,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 }));  // ../RTL/cortexm0ds_logic.v(20214)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100010011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1446|_al_u5927  (
    .a({open_n5244,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 }),
    .b({open_n5245,_al_u5926_o}),
    .c({_al_u1348_o,_al_u1445_o}),
    .d({_al_u1445_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [18],_al_u5927_o}));
  // ../RTL/cortexm0ds_logic.v(18858)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1448|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyrax6_reg  (
    .a({open_n5266,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .b({_al_u1447_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] }),
    .mi({open_n5277,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({_al_u1448_o,_al_u1447_o}),
    .q({open_n5282,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] }));  // ../RTL/cortexm0ds_logic.v(18858)
  // ../RTL/cortexm0ds_logic.v(18886)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1450|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eitax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 }),
    .mi({open_n5293,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({_al_u1450_o,_al_u2213_o}),
    .q({open_n5298,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[19] }));  // ../RTL/cortexm0ds_logic.v(18886)
  // ../RTL/cortexm0ds_logic.v(18783)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1452|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntnax6_reg  (
    .a({open_n5299,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1450_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1451_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1449_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] }),
    .mi({open_n5310,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({_al_u1452_o,_al_u1451_o}),
    .q({open_n5315,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] }));  // ../RTL/cortexm0ds_logic.v(18783)
  // ../RTL/cortexm0ds_logic.v(20233)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1453|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6_reg  (
    .a({_al_u1452_o,open_n5316}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ,_al_u4073_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 ,_al_u4071_o}),
    .f({_al_u1453_o,open_n5335}),
    .q({open_n5339,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 }));  // ../RTL/cortexm0ds_logic.v(20233)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(D*~C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100010011001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100010011001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1454|_al_u5938  (
    .a({open_n5340,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 }),
    .b({open_n5341,_al_u5937_o}),
    .c({_al_u1348_o,_al_u1453_o}),
    .d({_al_u1453_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [19],_al_u5938_o}));
  // ../RTL/cortexm0ds_logic.v(18885)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1455|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egtax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 }),
    .mi({open_n5369,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .f({_al_u1455_o,_al_u2221_o}),
    .q({open_n5385,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[20] }));  // ../RTL/cortexm0ds_logic.v(18885)
  // ../RTL/cortexm0ds_logic.v(17229)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~D)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(C*B*~D)"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1456|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X4jpw6_reg  (
    .b({_al_u1455_o,_al_u6926_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,_al_u6844_o}),
    .f({_al_u1456_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .q({open_n5408,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] }));  // ../RTL/cortexm0ds_logic.v(17229)
  // ../RTL/cortexm0ds_logic.v(17918)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1457|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T80qw6_reg  (
    .a({open_n5409,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1456_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[18] }),
    .mi({open_n5420,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .f({_al_u1457_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqyow6 }),
    .q({open_n5425,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[18] }));  // ../RTL/cortexm0ds_logic.v(17918)
  // ../RTL/cortexm0ds_logic.v(17228)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1460|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2jpw6_reg  (
    .a({open_n5426,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1458_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1459_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1457_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] }),
    .mi({open_n5437,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .f({_al_u1460_o,_al_u1459_o}),
    .q({open_n5442,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] }));  // ../RTL/cortexm0ds_logic.v(17228)
  // ../RTL/cortexm0ds_logic.v(19976)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1461|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6_reg  (
    .a({_al_u1460_o,open_n5443}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ,_al_u4078_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 ,_al_u4076_o}),
    .f({_al_u1461_o,open_n5462}),
    .q({open_n5466,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 }));  // ../RTL/cortexm0ds_logic.v(19976)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(D*~C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100010011001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100010011001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1462|_al_u5943  (
    .a({open_n5467,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 }),
    .b({open_n5468,_al_u5942_o}),
    .c({_al_u1348_o,_al_u1461_o}),
    .d({_al_u1461_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [20],_al_u5943_o}));
  // ../RTL/cortexm0ds_logic.v(18781)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1463|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npnax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] }),
    .mi({open_n5496,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .f({_al_u1463_o,_al_u2229_o}),
    .q({open_n5512,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[21] }));  // ../RTL/cortexm0ds_logic.v(18781)
  // ../RTL/cortexm0ds_logic.v(17298)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1465|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfkpw6_reg  (
    .a({open_n5513,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1464_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] }),
    .mi({open_n5524,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .f({_al_u1465_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhyow6 }),
    .q({open_n5529,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[19] }));  // ../RTL/cortexm0ds_logic.v(17298)
  // ../RTL/cortexm0ds_logic.v(18884)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1467|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eetax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 }),
    .mi({open_n5533,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .f({_al_u1467_o,_al_u2231_o}),
    .q({open_n5549,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[21] }));  // ../RTL/cortexm0ds_logic.v(18884)
  // ../RTL/cortexm0ds_logic.v(17528)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1468|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxopw6_reg  (
    .a({open_n5550,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1466_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1467_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1465_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] }),
    .mi({open_n5554,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .f({_al_u1468_o,_al_u1466_o}),
    .q({open_n5570,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[21] }));  // ../RTL/cortexm0ds_logic.v(17528)
  // ../RTL/cortexm0ds_logic.v(19986)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1469|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6_reg  (
    .a({_al_u1468_o,open_n5571}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ,_al_u4083_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ,_al_u4081_o}),
    .f({_al_u1469_o,open_n5586}),
    .q({open_n5590,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 }));  // ../RTL/cortexm0ds_logic.v(19986)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100010011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1470|_al_u5948  (
    .a({open_n5591,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 }),
    .b({open_n5592,_al_u5947_o}),
    .c({_al_u1348_o,_al_u1469_o}),
    .d({_al_u1469_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [21],_al_u5948_o}));
  // ../RTL/cortexm0ds_logic.v(20004)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1471|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1fbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] }),
    .mi({open_n5616,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u1471_o,_al_u2240_o}),
    .q({open_n5632,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[22] }));  // ../RTL/cortexm0ds_logic.v(20004)
  // ../RTL/cortexm0ds_logic.v(20011)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1472|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tffbx6_reg  (
    .a({open_n5633,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({_al_u1471_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] }),
    .mi({open_n5637,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u1472_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7yow6 }),
    .q({open_n5653,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[20] }));  // ../RTL/cortexm0ds_logic.v(20011)
  // ../RTL/cortexm0ds_logic.v(20010)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1476|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdfbx6_reg  (
    .a({open_n5654,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1474_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .c({_al_u1475_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] }),
    .mi({open_n5658,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u1476_o,_al_u1475_o}),
    .q({open_n5674,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[22] }));  // ../RTL/cortexm0ds_logic.v(20010)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1477|_al_u788  (
    .a({_al_u1476_o,open_n5675}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ,open_n5676}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1477_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [22]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(D*~C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100010011001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100010011001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1478|_al_u6208  (
    .a({open_n5701,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 }),
    .b({open_n5702,_al_u6207_o}),
    .c({_al_u1348_o,_al_u1477_o}),
    .d({_al_u1477_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [22],_al_u6208_o}));
  // ../RTL/cortexm0ds_logic.v(18768)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1479|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szmax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 }),
    .mi({open_n5730,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u1479_o,_al_u2248_o}),
    .q({open_n5746,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[23] }));  // ../RTL/cortexm0ds_logic.v(18768)
  // ../RTL/cortexm0ds_logic.v(18064)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1480|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gp6ax6_reg  (
    .b({_al_u1479_o,open_n5749}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,_al_u3769_o}),
    .mi({open_n5753,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u1480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 }),
    .q({open_n5769,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] }));  // ../RTL/cortexm0ds_logic.v(18064)
  // ../RTL/cortexm0ds_logic.v(18065)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1481|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr6ax6_reg  (
    .a({open_n5770,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[21] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] }),
    .mi({open_n5774,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u1481_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxow6 }),
    .q({open_n5790,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[21] }));  // ../RTL/cortexm0ds_logic.v(18065)
  // ../RTL/cortexm0ds_logic.v(18850)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1484|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qirax6_reg  (
    .a({open_n5791,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C96pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .c({_al_u1483_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1481_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] }),
    .mi({open_n5795,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u1484_o,_al_u1483_o}),
    .q({open_n5811,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] }));  // ../RTL/cortexm0ds_logic.v(18850)
  // ../RTL/cortexm0ds_logic.v(20096)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1485|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6_reg  (
    .a({_al_u1484_o,open_n5812}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ,_al_u4093_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 ,_al_u4091_o}),
    .f({_al_u1485_o,open_n5831}),
    .q({open_n5835,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 }));  // ../RTL/cortexm0ds_logic.v(20096)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100010011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1486|_al_u6198  (
    .a({open_n5836,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23]}),
    .b({open_n5837,_al_u6197_o}),
    .c({_al_u1348_o,_al_u1485_o}),
    .d({_al_u1485_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [23],_al_u6198_o}));
  // ../RTL/cortexm0ds_logic.v(18748)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1488|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvlax6_reg  (
    .a({open_n5858,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1487_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] }),
    .mi({open_n5869,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u1488_o,_al_u1487_o}),
    .q({open_n5874,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] }));  // ../RTL/cortexm0ds_logic.v(18748)
  // ../RTL/cortexm0ds_logic.v(17912)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1489|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Twzpw6_reg  (
    .a({open_n5875,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1488_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] }),
    .mi({open_n5886,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u1489_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voxow6 }),
    .q({open_n5891,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[22] }));  // ../RTL/cortexm0ds_logic.v(17912)
  // ../RTL/cortexm0ds_logic.v(18878)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1490|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2tax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 }),
    .mi({open_n5902,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u1490_o,_al_u2433_o}),
    .q({open_n5907,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[24] }));  // ../RTL/cortexm0ds_logic.v(18878)
  // ../RTL/cortexm0ds_logic.v(17665)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1492|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxspw6_reg  (
    .a({open_n5908,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .b({_al_u1490_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1491_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1489_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] }),
    .mi({open_n5919,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u1492_o,_al_u1491_o}),
    .q({open_n5924,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] }));  // ../RTL/cortexm0ds_logic.v(17665)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"))
    \_al_u1493|_al_u800  (
    .a({_al_u1492_o,open_n5925}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ,open_n5926}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1493_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [24]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1494|_al_u1601  (
    .c({_al_u1348_o,_al_u1348_o}),
    .d({_al_u1493_o,_al_u1600_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [24],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [5]}));
  // ../RTL/cortexm0ds_logic.v(18780)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1495|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnnax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] }),
    .mi({open_n5974,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u1495_o,_al_u2255_o}),
    .q({open_n5990,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[25] }));  // ../RTL/cortexm0ds_logic.v(18780)
  // ../RTL/cortexm0ds_logic.v(17916)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1496|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T40qw6_reg  (
    .a({open_n5991,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({_al_u1495_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] }),
    .mi({open_n5995,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u1496_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xow6 }),
    .q({open_n6011,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[23] }));  // ../RTL/cortexm0ds_logic.v(17916)
  // ../RTL/cortexm0ds_logic.v(17677)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1497|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbtpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,open_n6014}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] ,_al_u5871_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1496_o,_al_u7105_o}),
    .f({_al_u1497_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .q({open_n6035,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[23] }));  // ../RTL/cortexm0ds_logic.v(17677)
  // ../RTL/cortexm0ds_logic.v(18753)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1500|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5max6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .b({_al_u1497_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({_al_u1498_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1499_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] }),
    .mi({open_n6046,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u1500_o,_al_u1499_o}),
    .q({open_n6051,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] }));  // ../RTL/cortexm0ds_logic.v(18753)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100111100000011),
    .MODE("LOGIC"))
    \_al_u1501|_al_u2257  (
    .a({open_n6052,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] }),
    .d({_al_u1500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ,_al_u2257_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u1502|_al_u1593  (
    .c({_al_u1348_o,_al_u1348_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv ,_al_u1592_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [25],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [3]}));
  // ../RTL/cortexm0ds_logic.v(18749)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1504|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxlax6_reg  (
    .a({open_n6097,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1503_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] }),
    .mi({open_n6101,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u1504_o,_al_u1503_o}),
    .q({open_n6117,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] }));  // ../RTL/cortexm0ds_logic.v(18749)
  // ../RTL/cortexm0ds_logic.v(17913)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1505|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyzpw6_reg  (
    .a({open_n6118,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] }),
    .mi({open_n6129,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u1505_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynwow6 }),
    .q({open_n6134,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[24] }));  // ../RTL/cortexm0ds_logic.v(17913)
  // ../RTL/cortexm0ds_logic.v(18879)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1507|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4tax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 }),
    .mi({open_n6138,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u1507_o,_al_u2451_o}),
    .q({open_n6154,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[26] }));  // ../RTL/cortexm0ds_logic.v(18879)
  // ../RTL/cortexm0ds_logic.v(17693)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1508|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxtpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1505_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1507_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] }),
    .mi({open_n6158,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u1508_o,_al_u1506_o}),
    .q({open_n6174,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] }));  // ../RTL/cortexm0ds_logic.v(17693)
  // ../RTL/cortexm0ds_logic.v(19946)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b1100111100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1509|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6_reg  (
    .b({_al_u1334_o,_al_u4098_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1508_o,_al_u4096_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ,open_n6191}),
    .q({open_n6195,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 }));  // ../RTL/cortexm0ds_logic.v(19946)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1510|_al_u1574  (
    .c({_al_u1348_o,_al_u1348_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv ,_al_u1573_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [26],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [4]}));
  // ../RTL/cortexm0ds_logic.v(18880)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1511|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6tax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 }),
    .mi({open_n6234,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u1511_o,_al_u2441_o}),
    .q({open_n6239,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[27] }));  // ../RTL/cortexm0ds_logic.v(18880)
  // ../RTL/cortexm0ds_logic.v(17902)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1512|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zczpw6_reg  (
    .b({_al_u1511_o,_al_u7113_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] ,_al_u5906_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,_al_u7092_o}),
    .f({_al_u1512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .q({open_n6258,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] }));  // ../RTL/cortexm0ds_logic.v(17902)
  // ../RTL/cortexm0ds_logic.v(17914)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1513|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T00qw6_reg  (
    .a({open_n6259,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[25] }),
    .mi({open_n6270,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u1513_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdwow6 }),
    .q({open_n6275,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[25] }));  // ../RTL/cortexm0ds_logic.v(17914)
  // ../RTL/cortexm0ds_logic.v(18750)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1516|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xzlax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .b({_al_u1513_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({_al_u1514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1515_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] }),
    .mi({open_n6279,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u1516_o,_al_u1515_o}),
    .q({open_n6295,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] }));  // ../RTL/cortexm0ds_logic.v(18750)
  // ../RTL/cortexm0ds_logic.v(19941)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b1100111100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1517|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6_reg  (
    .b({_al_u1334_o,_al_u4103_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1516_o,_al_u4101_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ,open_n6312}),
    .q({open_n6316,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 }));  // ../RTL/cortexm0ds_logic.v(19941)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1518|_al_u1542  (
    .c({_al_u1348_o,_al_u1348_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv ,_al_u1541_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [27],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [30]}));
  // ../RTL/cortexm0ds_logic.v(20189)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1521|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pejbx6_reg  (
    .a({open_n6345,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] }),
    .mi({open_n6349,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({_al_u1521_o,_al_u2417_o}),
    .q({open_n6365,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[26] }));  // ../RTL/cortexm0ds_logic.v(20189)
  // ../RTL/cortexm0ds_logic.v(20170)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1522|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] }),
    .mi({open_n6376,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({_al_u1522_o,_al_u2416_o}),
    .q({open_n6381,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[28] }));  // ../RTL/cortexm0ds_logic.v(20170)
  // ../RTL/cortexm0ds_logic.v(20176)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1523|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rpibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] }),
    .mi({open_n6392,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({_al_u1523_o,_al_u2414_o}),
    .q({open_n6397,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[28] }));  // ../RTL/cortexm0ds_logic.v(20176)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1524|_al_u1536  (
    .b({_al_u1522_o,_al_u1535_o}),
    .c({_al_u1523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] }),
    .d({_al_u1521_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 }),
    .f({_al_u1524_o,_al_u1536_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"))
    \_al_u1525|_al_u824  (
    .a({_al_u1524_o,open_n6420}),
    .b({_al_u823_o,open_n6421}),
    .c({_al_u1334_o,_al_u823_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1525_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [28]}));
  // ../RTL/cortexm0ds_logic.v(17248)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1527|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmjpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 }),
    .mi({open_n6445,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u1527_o,_al_u2425_o}),
    .q({open_n6461,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[29] }));  // ../RTL/cortexm0ds_logic.v(17248)
  // ../RTL/cortexm0ds_logic.v(17903)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1528|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zezpw6_reg  (
    .b({_al_u1527_o,_al_u7097_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] ,_al_u5866_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,_al_u7092_o}),
    .f({_al_u1528_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .q({open_n6480,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] }));  // ../RTL/cortexm0ds_logic.v(17903)
  // ../RTL/cortexm0ds_logic.v(17915)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1529|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T20qw6_reg  (
    .a({open_n6481,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1528_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[27] }),
    .mi({open_n6485,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u1529_o,_al_u2427_o}),
    .q({open_n6501,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[27] }));  // ../RTL/cortexm0ds_logic.v(17915)
  // ../RTL/cortexm0ds_logic.v(18751)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1532|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1max6_reg  (
    .a({open_n6502,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eq4pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({_al_u1531_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1529_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] }),
    .mi({open_n6506,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u1532_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eq4pw6 }),
    .q({open_n6522,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] }));  // ../RTL/cortexm0ds_logic.v(18751)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"))
    \_al_u1533|_al_u830  (
    .a({_al_u1532_o,open_n6523}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ,open_n6524}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1533_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [29]}));
  // ../RTL/cortexm0ds_logic.v(18741)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1535|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cilax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] }),
    .mi({open_n6548,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({_al_u1535_o,_al_u2268_o}),
    .q({open_n6564,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[30] }));  // ../RTL/cortexm0ds_logic.v(18741)
  // ../RTL/cortexm0ds_logic.v(17894)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1537|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Exypw6_reg  (
    .a({open_n6565,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1536_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] }),
    .mi({open_n6569,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({_al_u1537_o,_al_u2267_o}),
    .q({open_n6585,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[28] }));  // ../RTL/cortexm0ds_logic.v(17894)
  // ../RTL/cortexm0ds_logic.v(17216)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1540|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoipw6_reg  (
    .a({open_n6586,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1538_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1539_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1537_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] }),
    .mi({open_n6597,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({_al_u1540_o,_al_u1539_o}),
    .q({open_n6602,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] }));  // ../RTL/cortexm0ds_logic.v(17216)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1541|_al_u836  (
    .a({_al_u1540_o,open_n6603}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ,open_n6604}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1541_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [30]}));
  // ../RTL/cortexm0ds_logic.v(18876)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1543|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hysax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] }),
    .mi({open_n6639,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1543_o,_al_u1946_o}),
    .q({open_n6644,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[6] }));  // ../RTL/cortexm0ds_logic.v(18876)
  // ../RTL/cortexm0ds_logic.v(17898)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1545|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B5zpw6_reg  (
    .a({open_n6645,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1544_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] }),
    .mi({open_n6649,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1545_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq0pw6 }),
    .q({open_n6665,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[4] }));  // ../RTL/cortexm0ds_logic.v(17898)
  // ../RTL/cortexm0ds_logic.v(17640)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1548|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3spw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1545_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .c({_al_u1546_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1547_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] }),
    .mi({open_n6669,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1548_o,_al_u1546_o}),
    .q({open_n6685,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[6] }));  // ../RTL/cortexm0ds_logic.v(17640)
  // ../RTL/cortexm0ds_logic.v(19812)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b1100111100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1549|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6_reg  (
    .b({_al_u1334_o,_al_u4143_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1548_o,_al_u4141_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ,open_n6702}),
    .q({open_n6706,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 }));  // ../RTL/cortexm0ds_logic.v(19812)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*C*A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0100110011001100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u1550|_al_u5891  (
    .a({open_n6707,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 }),
    .b({open_n6708,_al_u5890_o}),
    .c({_al_u1348_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [6],_al_u5891_o}));
  // ../RTL/cortexm0ds_logic.v(20180)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1551|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] }),
    .mi({open_n6732,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({_al_u1551_o,_al_u1974_o}),
    .q({open_n6748,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[9] }));  // ../RTL/cortexm0ds_logic.v(20180)
  // ../RTL/cortexm0ds_logic.v(20182)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1553|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1jbx6_reg  (
    .a({open_n6749,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1552_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] }),
    .mi({open_n6753,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({_al_u1553_o,_al_u1975_o}),
    .q({open_n6769,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[7] }));  // ../RTL/cortexm0ds_logic.v(20182)
  // ../RTL/cortexm0ds_logic.v(17947)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1554|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ht1qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 }),
    .mi({open_n6773,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({_al_u1554_o,_al_u1972_o}),
    .q({open_n6789,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[9] }));  // ../RTL/cortexm0ds_logic.v(17947)
  // ../RTL/cortexm0ds_logic.v(20179)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1556|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .b({_al_u1553_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({_al_u1554_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1555_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] }),
    .mi({open_n6800,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({_al_u1556_o,_al_u1555_o}),
    .q({open_n6805,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[9] }));  // ../RTL/cortexm0ds_logic.v(20179)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100111100000011),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u1558|_al_u1557  (
    .b({open_n6808,_al_u1334_o}),
    .c({_al_u1348_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ,_al_u1556_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(18852)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1560|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmrax6_reg  (
    .a({open_n6829,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .b({_al_u1559_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] }),
    .mi({open_n6840,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u1560_o,_al_u1559_o}),
    .q({open_n6845,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] }));  // ../RTL/cortexm0ds_logic.v(18852)
  // ../RTL/cortexm0ds_logic.v(17893)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1561|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evypw6_reg  (
    .a({open_n6846,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1560_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] }),
    .mi({open_n6857,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u1561_o,_al_u2279_o}),
    .q({open_n6862,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[29] }));  // ../RTL/cortexm0ds_logic.v(17893)
  // ../RTL/cortexm0ds_logic.v(17523)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1562|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnopw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] }),
    .mi({open_n6873,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u1562_o,_al_u2277_o}),
    .q({open_n6878,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[31] }));  // ../RTL/cortexm0ds_logic.v(17523)
  // ../RTL/cortexm0ds_logic.v(17455)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1564|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efnpw6_reg  (
    .a({open_n6879,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1562_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1563_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1561_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] }),
    .mi({open_n6883,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u1564_o,_al_u1563_o}),
    .q({open_n6899,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] }));  // ../RTL/cortexm0ds_logic.v(17455)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1565|_al_u854  (
    .a({_al_u1564_o,open_n6900}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ,open_n6901}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [31]}));
  // ../RTL/cortexm0ds_logic.v(18767)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1568|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Txmax6_reg  (
    .a({open_n6926,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({_al_u1567_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] }),
    .mi({open_n6937,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1568_o,_al_u1567_o}),
    .q({open_n6942,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] }));  // ../RTL/cortexm0ds_logic.v(18767)
  // ../RTL/cortexm0ds_logic.v(17895)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1569|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezypw6_reg  (
    .a({open_n6943,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1568_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] }),
    .mi({open_n6947,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1569_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kp1pw6 }),
    .q({open_n6963,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[2] }));  // ../RTL/cortexm0ds_logic.v(17895)
  // ../RTL/cortexm0ds_logic.v(18869)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1571|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lksax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 }),
    .mi({open_n6974,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1571_o,_al_u1928_o}),
    .q({open_n6979,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[4] }));  // ../RTL/cortexm0ds_logic.v(18869)
  // ../RTL/cortexm0ds_logic.v(17224)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1572|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuipw6_reg  (
    .a({open_n6980,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1570_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({_al_u1571_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1569_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] }),
    .mi({open_n6991,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1572_o,_al_u1570_o}),
    .q({open_n6996,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] }));  // ../RTL/cortexm0ds_logic.v(17224)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"))
    \_al_u1573|_al_u860  (
    .a({_al_u1572_o,open_n6997}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ,open_n6998}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1573_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [4]}));
  // ../RTL/cortexm0ds_logic.v(18766)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1575|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvmax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] }),
    .mi({open_n7029,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u1575_o,_al_u1910_o}),
    .q({open_n7034,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[2] }));  // ../RTL/cortexm0ds_logic.v(18766)
  // ../RTL/cortexm0ds_logic.v(17904)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1576|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgzpw6_reg  (
    .b({_al_u1575_o,open_n7037}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,_al_u7032_o}),
    .f({_al_u1576_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .q({open_n7058,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] }));  // ../RTL/cortexm0ds_logic.v(17904)
  // ../RTL/cortexm0ds_logic.v(17892)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1577|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftypw6_reg  (
    .a({open_n7059,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1576_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[0] }),
    .mi({open_n7070,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u1577_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro2pw6 }),
    .q({open_n7075,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[0] }));  // ../RTL/cortexm0ds_logic.v(17892)
  // ../RTL/cortexm0ds_logic.v(17684)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1580|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yftpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1577_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .c({_al_u1578_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1579_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] }),
    .mi({open_n7079,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u1580_o,_al_u1578_o}),
    .q({open_n7095,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[2] }));  // ../RTL/cortexm0ds_logic.v(17684)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1584|_al_u1583  (
    .b({_al_u1583_o,open_n7098}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u1582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u1584_o,_al_u1583_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b1100111100000011),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u1585|_al_u1581  (
    .b({_al_u1348_o,_al_u1334_o}),
    .c({_al_u1584_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 }),
    .d({_al_u1581_o,_al_u1580_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [2],_al_u1581_o}));
  // ../RTL/cortexm0ds_logic.v(17896)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1588|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1zpw6_reg  (
    .a({open_n7141,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1587_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] }),
    .mi({open_n7152,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1588_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X62pw6 }),
    .q({open_n7157,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[1] }));  // ../RTL/cortexm0ds_logic.v(17896)
  // ../RTL/cortexm0ds_logic.v(17420)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1589|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbmpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] }),
    .mi({open_n7168,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1589_o,_al_u1921_o}),
    .q({open_n7173,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[3] }));  // ../RTL/cortexm0ds_logic.v(17420)
  // ../RTL/cortexm0ds_logic.v(17421)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1591|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdmpw6_reg  (
    .a({open_n7174,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .b({_al_u1589_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .c({_al_u1590_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1588_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] }),
    .mi({open_n7185,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1591_o,_al_u1590_o}),
    .q({open_n7190,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] }));  // ../RTL/cortexm0ds_logic.v(17421)
  // ../RTL/cortexm0ds_logic.v(18874)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1592|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jusax6_reg  (
    .a({_al_u1591_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 }),
    .mi({open_n7201,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1592_o,_al_u1919_o}),
    .q({open_n7206,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[3] }));  // ../RTL/cortexm0ds_logic.v(18874)
  // ../RTL/cortexm0ds_logic.v(17897)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1596|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3zpw6_reg  (
    .a({open_n7207,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1595_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] }),
    .mi({open_n7211,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1596_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X71pw6 }),
    .q({open_n7227,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[3] }));  // ../RTL/cortexm0ds_logic.v(17897)
  // ../RTL/cortexm0ds_logic.v(18773)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1598|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9nax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] }),
    .mi({open_n7238,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1598_o,_al_u1939_o}),
    .q({open_n7243,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[5] }));  // ../RTL/cortexm0ds_logic.v(18773)
  // ../RTL/cortexm0ds_logic.v(17525)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1599|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Propw6_reg  (
    .a({open_n7244,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1597_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .c({_al_u1598_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1596_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] }),
    .mi({open_n7248,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1599_o,_al_u1597_o}),
    .q({open_n7264,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] }));  // ../RTL/cortexm0ds_logic.v(17525)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1600|_al_u878  (
    .a({_al_u1599_o,open_n7265}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ,open_n7266}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1600_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [5]}));
  // ../RTL/cortexm0ds_logic.v(17934)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1604|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O41qw6_reg  (
    .a({open_n7291,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1603_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] }),
    .mi({open_n7295,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({_al_u1604_o,_al_u1899_o}),
    .q({open_n7311,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[6] }));  // ../RTL/cortexm0ds_logic.v(17934)
  // ../RTL/cortexm0ds_logic.v(17931)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1605|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry0qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] }),
    .mi({open_n7315,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({_al_u1605_o,_al_u1893_o}),
    .q({open_n7331,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[8] }));  // ../RTL/cortexm0ds_logic.v(17931)
  // ../RTL/cortexm0ds_logic.v(18894)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1606|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eytax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 }),
    .mi({open_n7342,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({_al_u1606_o,_al_u1895_o}),
    .q({open_n7347,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[8] }));  // ../RTL/cortexm0ds_logic.v(18894)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1607|_al_u2288  (
    .a({open_n7348,_al_u2284_o}),
    .b({_al_u1605_o,_al_u2285_o}),
    .c({_al_u1606_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peqow6 }),
    .d({_al_u1604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ciqow6 }),
    .f({_al_u1607_o,_al_u2288_o}));
  // ../RTL/cortexm0ds_logic.v(17935)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1608|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6_reg  (
    .a({_al_u1607_o,open_n7373}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ,_al_u4108_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ,_al_u4106_o}),
    .f({_al_u1608_o,open_n7388}),
    .q({open_n7392,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 }));  // ../RTL/cortexm0ds_logic.v(17935)
  // ../RTL/cortexm0ds_logic.v(17911)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1611|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uuzpw6_reg  (
    .a({open_n7393,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({_al_u1610_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] }),
    .mi({open_n7397,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u1611_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80pw6 }),
    .q({open_n7413,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[5] }));  // ../RTL/cortexm0ds_logic.v(17911)
  // ../RTL/cortexm0ds_logic.v(17899)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1612|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A7zpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,open_n7416}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1611_o,_al_u3769_o}),
    .mi({open_n7427,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u1612_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 }),
    .q({open_n7432,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[5] }));  // ../RTL/cortexm0ds_logic.v(17899)
  // ../RTL/cortexm0ds_logic.v(17629)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1614|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bsrpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] }),
    .mi({open_n7436,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u1614_o,_al_u1957_o}),
    .q({open_n7452,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[7] }));  // ../RTL/cortexm0ds_logic.v(17629)
  // ../RTL/cortexm0ds_logic.v(18877)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1615|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0tax6_reg  (
    .a({open_n7453,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({_al_u1613_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .c({_al_u1614_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1612_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] }),
    .mi({open_n7457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u1615_o,_al_u1613_o}),
    .q({open_n7473,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] }));  // ../RTL/cortexm0ds_logic.v(18877)
  // ../RTL/cortexm0ds_logic.v(17718)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1616|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6_reg  (
    .a({_al_u1615_o,open_n7474}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ,_al_u4123_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ,_al_u4121_o}),
    .f({_al_u1616_o,open_n7493}),
    .q({open_n7497,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 }));  // ../RTL/cortexm0ds_logic.v(17718)
  // ../RTL/cortexm0ds_logic.v(17852)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1618|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqxpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] }),
    .mi({open_n7508,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({_al_u1618_o,_al_u2033_o}),
    .q({open_n7513,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[10] }));  // ../RTL/cortexm0ds_logic.v(17852)
  // ../RTL/cortexm0ds_logic.v(17854)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1620|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Huxpw6_reg  (
    .a({open_n7514,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1619_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] }),
    .mi({open_n7518,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({_al_u1620_o,_al_u2037_o}),
    .q({open_n7534,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[8] }));  // ../RTL/cortexm0ds_logic.v(17854)
  // ../RTL/cortexm0ds_logic.v(18790)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1621|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7oax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] }),
    .mi({open_n7545,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({_al_u1621_o,_al_u2036_o}),
    .q({open_n7550,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[10] }));  // ../RTL/cortexm0ds_logic.v(18790)
  // ../RTL/cortexm0ds_logic.v(18865)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1623|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocsax6_reg  (
    .a({open_n7551,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .b({_al_u1621_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .c({_al_u1622_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1620_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] }),
    .mi({open_n7562,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({_al_u1623_o,_al_u1622_o}),
    .q({open_n7567,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[10] }));  // ../RTL/cortexm0ds_logic.v(18865)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0111111101110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0111111101110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1624|_al_u896  (
    .a({_al_u1623_o,open_n7568}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ,open_n7569}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1624_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [10]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*B*~A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~(D*B*~A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1011000011110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1011000011110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1625|_al_u6182  (
    .a({open_n7594,_al_u1624_o}),
    .b({open_n7595,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10]}),
    .c({_al_u1348_o,_al_u6181_o}),
    .d({_al_u1624_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [10],_al_u6182_o}));
  // ../RTL/cortexm0ds_logic.v(19801)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1626|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zp8bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] }),
    .mi({open_n7630,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .f({_al_u1626_o,_al_u2059_o}),
    .q({open_n7635,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[11] }));  // ../RTL/cortexm0ds_logic.v(19801)
  // ../RTL/cortexm0ds_logic.v(19802)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1627|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zr8bx6_reg  (
    .b({_al_u1626_o,_al_u6994_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] ,_al_u6188_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,_al_u6969_o}),
    .f({_al_u1627_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .q({open_n7654,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] }));  // ../RTL/cortexm0ds_logic.v(19802)
  // ../RTL/cortexm0ds_logic.v(19803)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1628|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt8bx6_reg  (
    .a({open_n7655,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1627_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[9] }),
    .mi({open_n7659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .f({_al_u1628_o,_al_u2060_o}),
    .q({open_n7675,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[9] }));  // ../RTL/cortexm0ds_logic.v(19803)
  // ../RTL/cortexm0ds_logic.v(19771)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1629|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc7bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] }),
    .mi({open_n7686,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .f({_al_u1629_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hy1pw6 }),
    .q({open_n7691,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[11] }));  // ../RTL/cortexm0ds_logic.v(19771)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1631|_al_u293  (
    .b({_al_u1629_o,open_n7694}),
    .c({_al_u1630_o,\u_cmsdk_mcu/u_ahb_rom/we }),
    .d({_al_u1628_o,\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [12]}),
    .f({_al_u1631_o,\u_cmsdk_mcu/u_ahb_rom/n16 }));
  // ../RTL/cortexm0ds_logic.v(19765)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(~D*~((B*A))*~(C)+~D*(B*A)*~(C)+~(~D)*(B*A)*C+~D*(B*A)*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0111111101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1632|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6_reg  (
    .a({_al_u1631_o,open_n7715}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ,_al_u4118_o}),
    .c({_al_u1334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ,_al_u4116_o}),
    .f({_al_u1632_o,open_n7730}),
    .q({open_n7734,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 }));  // ../RTL/cortexm0ds_logic.v(19765)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*B*~A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~(D*B*~A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1011000011110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1011000011110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1633|_al_u6187  (
    .a({open_n7735,_al_u1632_o}),
    .b({open_n7736,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 }),
    .c({_al_u1348_o,_al_u6186_o}),
    .d({_al_u1632_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [11],_al_u6187_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~(D*A)))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(C*~(~B*~(D*A)))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1110000011000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1636|_al_u1375  (
    .a({open_n7761,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u1636_o,_al_u1375_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(B*~(~D*C)))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~A*~(B*~(~D*C)))"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b0001000101010001),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0001000101010001),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1637|_al_u1634  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb1ju6 ,_al_u1363_o}),
    .b({_al_u1634_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({_al_u1635_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u1636_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ,_al_u1634_o}));
  // ../RTL/cortexm0ds_logic.v(18692)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1638|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6_reg  (
    .b({_al_u1359_o,_al_u1638_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Srbow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 }),
    .f({_al_u1638_o,open_n7825}),
    .q({open_n7829,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }));  // ../RTL/cortexm0ds_logic.v(18692)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u1640|_al_u1790  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17771)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1641|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 }),
    .q({open_n7873,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 }));  // ../RTL/cortexm0ds_logic.v(17771)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1642|_al_u7203  (
    .a({open_n7874,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [28]}),
    .f({_al_u1642_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfziu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(D*C*B*~A)"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0100000000000000),
    .MODE("LOGIC"))
    \_al_u1643|_al_u7171  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ,_al_u4289_o}),
    .b({_al_u1642_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [30]}),
    .f({_al_u1643_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ow6 }));
  // ../RTL/cortexm0ds_logic.v(17891)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(~A*~(~D*C)))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("~(B*~(~A*~(~D*C)))"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100110111),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0111011100110111),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1644|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6_reg  (
    .a({open_n7919,_al_u1644_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7aiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ,_al_u1648_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy9iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1643_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8aiu6_lutinv }),
    .f({_al_u1644_o,open_n7937}),
    .q({open_n7941,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 }));  // ../RTL/cortexm0ds_logic.v(17891)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~A*~(D*~C*B))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0101000101010101),
    .MODE("LOGIC"))
    \_al_u1647|_al_u1646  (
    .a({_al_u1646_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7aiu6_lutinv ,_al_u1646_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*~A))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~(C*B)*~(D*~A))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .INIT_LUTF0(16'b0010101000111111),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0010101000111111),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1652|_al_u1654  (
    .a({_al_u1360_o,_al_u1360_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb1ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .f({_al_u1652_o,_al_u1654_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1657|_al_u1656  (
    .a({open_n7986,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv }),
    .b({_al_u604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u1346_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u1656_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u1657_o,_al_u1656_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~D*~A*~(C*B))"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0000000000010101),
    .MODE("LOGIC"))
    \_al_u1661|_al_u1660  (
    .a({_al_u1659_o,open_n8011}),
    .b({_al_u679_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u1660_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ,_al_u1660_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(B*~A*~(~D*C))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0100010000000100),
    .MODE("LOGIC"))
    \_al_u1664|_al_u1663  (
    .a({_al_u1657_o,open_n8032}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u1663_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,_al_u1662_o}),
    .f({_al_u1664_o,_al_u1663_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~((~D*A))*~(C)+B*(~D*A)*~(C)+~(B)*(~D*A)*C+B*(~D*A)*C)"),
    //.LUTF1("(D*~(~A*~(C*~B)))"),
    //.LUTG0("~(B*~((~D*A))*~(C)+B*(~D*A)*~(C)+~(B)*(~D*A)*C+B*(~D*A)*C)"),
    //.LUTG1("(D*~(~A*~(C*~B)))"),
    .INIT_LUTF0(16'b1111001101010011),
    .INIT_LUTF1(16'b1011101000000000),
    .INIT_LUTG0(16'b1111001101010011),
    .INIT_LUTG1(16'b1011101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1668|_al_u1667  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv }),
    .b({_al_u1667_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u1668_o,_al_u1667_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B*A))"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(D*~(C*~B*A))"),
    //.LUTG1("(C*~(~B*D))"),
    .INIT_LUTF0(16'b1101111100000000),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b1101111100000000),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1669|_al_u3022  (
    .a({open_n8077,_al_u2461_o}),
    .b({_al_u1668_o,_al_u3015_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,_al_u3021_o}),
    .d({_al_u1664_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqfhu6 ,_al_u3022_o}));
  // ../RTL/cortexm0ds_logic.v(17587)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1670|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6_reg  (
    .a({open_n8102,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 }),
    .mi({open_n8114,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u1670_o,_al_u2470_o}),
    .q({open_n8118,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6 }));  // ../RTL/cortexm0ds_logic.v(17587)
  // ../RTL/cortexm0ds_logic.v(18361)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*C*~A))"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110011001100),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1671|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6_reg  (
    .a({_al_u1253_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 }),
    .b({_al_u1670_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 ,open_n8132}),
    .q({open_n8136,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 }));  // ../RTL/cortexm0ds_logic.v(18361)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1673|_al_u1254  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~(~C*B)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(A*~(D*~(~C*B)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000100010101010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000100010101010),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1674|_al_u2468  (
    .a({open_n8165,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv }),
    .b({open_n8166,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yn3iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 }),
    .d({_al_u1253_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ,_al_u2468_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1675|_al_u1731  (
    .b({open_n8193,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 }),
    .f({_al_u1675_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 }));
  // ../RTL/cortexm0ds_logic.v(18015)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0010111000111111),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0010111000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1677|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6_reg  (
    .a({_al_u1253_o,open_n8218}),
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 }),
    .mi({open_n8222,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yg3iu6 ,_al_u3872_o}),
    .q({open_n8238,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6 }));  // ../RTL/cortexm0ds_logic.v(18015)
  // ../RTL/cortexm0ds_logic.v(18008)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b0010001111101111),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b0010001111101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1679|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6_reg  (
    .a({_al_u1253_o,open_n8239}),
    .b({_al_u1676_o,_al_u1679_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .f({_al_u1679_o,open_n8258}),
    .q({open_n8262,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bx2qw6 }));  // ../RTL/cortexm0ds_logic.v(18008)
  // ../RTL/cortexm0ds_logic.v(17187)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1682|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6_reg  (
    .a({open_n8263,_al_u1826_o}),
    .b({open_n8264,_al_u1827_o}),
    .c({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1253_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,open_n8279}),
    .q({open_n8283,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 }));  // ../RTL/cortexm0ds_logic.v(17187)
  // ../RTL/cortexm0ds_logic.v(17938)
  EG_PHY_MSLICE #(
    //.LUT0("(D*A*~(~C*~B))"),
    //.LUT1("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000000000),
    .INIT_LUT1(16'b0010001111101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1685|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6_reg  (
    .a({_al_u1253_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 }),
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .mi({open_n8294,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 }),
    .f({_al_u1685_o,_al_u4025_o}),
    .q({open_n8299,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6 }));  // ../RTL/cortexm0ds_logic.v(17938)
  // ../RTL/cortexm0ds_logic.v(17188)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1689|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6_reg  (
    .b({_al_u1676_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,_al_u1675_o}),
    .mi({open_n8305,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W6ipw6 }),
    .f({_al_u1689_o,_al_u1823_o}),
    .q({open_n8321,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 }));  // ../RTL/cortexm0ds_logic.v(17188)
  // ../RTL/cortexm0ds_logic.v(18123)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001111101111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0010001111101111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1694|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6_reg  (
    .a({open_n8322,_al_u1253_o}),
    .b({_al_u1676_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 }),
    .mi({open_n8326,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 }),
    .f({_al_u1694_o,_al_u1697_o}),
    .q({open_n8342,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6 }));  // ../RTL/cortexm0ds_logic.v(18123)
  // ../RTL/cortexm0ds_logic.v(19932)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010111000111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1703|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6_reg  (
    .a({open_n8343,_al_u1253_o}),
    .b({_al_u1676_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 }),
    .mi({open_n8354,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 }),
    .f({_al_u1703_o,_al_u1706_o}),
    .q({open_n8359,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6 }));  // ../RTL/cortexm0ds_logic.v(19932)
  // ../RTL/cortexm0ds_logic.v(19985)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1712|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6_reg  (
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,_al_u1715_o}),
    .mi({open_n8365,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 }),
    .f({_al_u1712_o,_al_u1716_o}),
    .q({open_n8381,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 }));  // ../RTL/cortexm0ds_logic.v(19985)
  // ../RTL/cortexm0ds_logic.v(18099)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~B*~(D*A))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111001111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1715|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6_reg  (
    .a({open_n8382,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .b({_al_u1676_o,_al_u1675_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yg3iu6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 }),
    .f({_al_u1715_o,open_n8397}),
    .q({open_n8401,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 }));  // ../RTL/cortexm0ds_logic.v(18099)
  // ../RTL/cortexm0ds_logic.v(17310)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1720|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6_reg  (
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,_al_u1724_o}),
    .f({_al_u1720_o,open_n8418}),
    .q({open_n8422,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 }));  // ../RTL/cortexm0ds_logic.v(17310)
  // ../RTL/cortexm0ds_logic.v(17999)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1723|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6_reg  (
    .a({open_n8423,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 }),
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 }),
    .mi({open_n8434,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 }),
    .f({_al_u1723_o,_al_u368_o}),
    .q({open_n8439,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6 }));  // ../RTL/cortexm0ds_logic.v(17999)
  // ../RTL/cortexm0ds_logic.v(19944)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1726|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6_reg  (
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,_al_u1730_o}),
    .f({_al_u1726_o,open_n8460}),
    .q({open_n8464,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 }));  // ../RTL/cortexm0ds_logic.v(19944)
  // ../RTL/cortexm0ds_logic.v(17998)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1727|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1726_o,_al_u1727_o}),
    .f({_al_u1727_o,open_n8481}),
    .q({open_n8485,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn2qw6 }));  // ../RTL/cortexm0ds_logic.v(17998)
  // ../RTL/cortexm0ds_logic.v(19959)
  EG_PHY_MSLICE #(
    //.LUT0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001111101111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1730|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6_reg  (
    .a({open_n8486,_al_u1253_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P92iu6 ,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 }),
    .mi({open_n8497,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u1730_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P92iu6 }),
    .q({open_n8501,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpcbx6 }));  // ../RTL/cortexm0ds_logic.v(19959)
  // ../RTL/cortexm0ds_logic.v(17555)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1733|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6_reg  (
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,_al_u1737_o}),
    .f({_al_u1733_o,open_n8522}),
    .q({open_n8526,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 }));  // ../RTL/cortexm0ds_logic.v(17555)
  // ../RTL/cortexm0ds_logic.v(19943)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1734|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1733_o,_al_u1734_o}),
    .f({_al_u1734_o,open_n8547}),
    .q({open_n8551,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 }));  // ../RTL/cortexm0ds_logic.v(19943)
  // ../RTL/cortexm0ds_logic.v(17596)
  EG_PHY_MSLICE #(
    //.LUT0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001111101111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1737|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6_reg  (
    .a({open_n8552,_al_u1253_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52iu6 ,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 }),
    .mi({open_n8563,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 }),
    .f({_al_u1737_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52iu6 }),
    .q({open_n8568,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6 }));  // ../RTL/cortexm0ds_logic.v(17596)
  // ../RTL/cortexm0ds_logic.v(18048)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010111000111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0010111000111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1741|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6_reg  (
    .a({open_n8569,_al_u1253_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P22iu6 ,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F42iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 }),
    .mi({open_n8573,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 }),
    .f({_al_u1741_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P22iu6 }),
    .q({open_n8589,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6 }));  // ../RTL/cortexm0ds_logic.v(18048)
  // ../RTL/cortexm0ds_logic.v(17404)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0010111000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0010111000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1748|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6_reg  (
    .a({_al_u1253_o,open_n8590}),
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ,_al_u1749_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tj1iu6 ,open_n8609}),
    .q({open_n8613,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 }));  // ../RTL/cortexm0ds_logic.v(17404)
  // ../RTL/cortexm0ds_logic.v(17969)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1749|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tj1iu6 ,open_n8616}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 }),
    .mi({open_n8627,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u1749_o,_al_u1743_o}),
    .q({open_n8631,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T82qw6 }));  // ../RTL/cortexm0ds_logic.v(17969)
  // ../RTL/cortexm0ds_logic.v(18357)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101110111011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1751|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,_al_u5103_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ,_al_u5308_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 }),
    .f({_al_u1751_o,open_n8646}),
    .q({open_n8650,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vefax6 }));  // ../RTL/cortexm0ds_logic.v(18357)
  // ../RTL/cortexm0ds_logic.v(17405)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUT1("(B*~(A*~(D*~C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010111000111111),
    .INIT_LUT1(16'b0100110001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1753|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93iu6 ,_al_u1253_o}),
    .b({_al_u1752_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 }),
    .mi({open_n8661,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 }),
    .f({_al_u1753_o,_al_u1752_o}),
    .q({open_n8666,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6 }));  // ../RTL/cortexm0ds_logic.v(17405)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1755|_al_u529  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .d({_al_u529_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .f({_al_u1755_o,_al_u529_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~C*(D@B)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~A*~(~C*(D@B)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0101010001010001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0101010001010001),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1756|_al_u2307  (
    .a({open_n8695,_al_u1253_o}),
    .b({open_n8696,_al_u1755_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ,_al_u1761_o}),
    .d({_al_u1755_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .f({_al_u1756_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Spyhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~A*~(D*C*B))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"))
    \_al_u1758|_al_u1757  (
    .a({_al_u1756_o,open_n8721}),
    .b({_al_u1757_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .f({_al_u1758_o,_al_u1757_o}));
  // ../RTL/cortexm0ds_logic.v(17362)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(~D*B)))"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("~(~A*~(C*~(~D*B)))"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101010111010),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1111101010111010),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1761|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ,_al_u4032_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u1761_o,open_n8759}),
    .q({open_n8763,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 }));  // ../RTL/cortexm0ds_logic.v(17362)
  // ../RTL/cortexm0ds_logic.v(17380)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(~B*(C@(D*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b0001001000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1762|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6_reg  (
    .a({_al_u1756_o,_al_u1759_o}),
    .b({_al_u1761_o,_al_u1762_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ,_al_u1763_o}),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u1762_o,open_n8777}),
    .q({open_n8781,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 }));  // ../RTL/cortexm0ds_logic.v(17380)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1763|_al_u1760  (
    .b({open_n8784,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 }),
    .f({_al_u1763_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cayhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1765|_al_u1766  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 }),
    .d({_al_u1383_o,_al_u1765_o}),
    .f({_al_u1765_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17215)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~(D*~A))"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("~(C*B*~(D*~A))"),
    //.LUTG1("(~A*~(D*C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111100111111),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b0111111100111111),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1767|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ,_al_u1767_o}),
    .b({_al_u916_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,_al_u1770_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv }),
    .f({_al_u1767_o,open_n8846}),
    .q({open_n8850,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 }));  // ../RTL/cortexm0ds_logic.v(17215)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1768|_al_u919  (
    .a({_al_u696_o,open_n8851}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .f({_al_u1768_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(A*~(B*~(D*~C)))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(A*~(B*~(D*~C)))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0010101000100010),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0010101000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1770|_al_u1769  (
    .a({_al_u1768_o,open_n8876}),
    .b({_al_u1769_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u1770_o,_al_u1769_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1774|_al_u1773  (
    .b({open_n8903,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 ,_al_u1772_o}),
    .f({_al_u1774_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1777|_al_u1775  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u1775_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .f({_al_u1777_o,_al_u1775_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1110101000000000),
    .MODE("LOGIC"))
    \_al_u1779|_al_u1778  (
    .a({_al_u1778_o,open_n8954}),
    .b({_al_u933_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ,_al_u1774_o}),
    .f({_al_u1779_o,_al_u1778_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1782|_al_u1781  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u1781_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u1782_o,_al_u1781_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*A*~(~D*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*A*~(~D*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1010000000100000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1783|_al_u3397  (
    .a({open_n8999,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 }),
    .b({open_n9000,_al_u1783_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ,_al_u3396_o}),
    .d({_al_u1782_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u1783_o,_al_u3397_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1784|_al_u3816  (
    .a({open_n9025,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .b({open_n9026,_al_u1783_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,_al_u2849_o}),
    .d({_al_u1783_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({_al_u1784_o,_al_u3816_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1787|_al_u1785  (
    .a({_al_u906_o,_al_u606_o}),
    .b({_al_u1785_o,_al_u607_o}),
    .c({_al_u932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u1787_o,_al_u1785_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*~(D*C*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*~(D*C*B))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0010101010101010),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1788|_al_u1776  (
    .a({_al_u1787_o,open_n9075}),
    .b({_al_u1775_o,open_n9076}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u1788_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u1789|_al_u6705  (
    .c({_al_u1788_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 }),
    .d({_al_u1784_o,_al_u1781_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("~((B*A)*~(C)*~(D)+(B*A)*C*~(D)+~((B*A))*C*D+(B*A)*C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("~((B*A)*~(C)*~(D)+(B*A)*C*~(D)+~((B*A))*C*D+(B*A)*C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000111101110111),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000111101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1792|_al_u4259  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ,open_n9125}),
    .b({_al_u1791_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bofiu6_lutinv ,_al_u4259_o}));
  // ../RTL/cortexm0ds_logic.v(20244)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1793|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ,_al_u1794_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bofiu6_lutinv ,_al_u1793_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1793_o,open_n9165}),
    .q({open_n9169,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 }));  // ../RTL/cortexm0ds_logic.v(20244)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1794|_al_u353  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,open_n9172}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg }),
    .d({_al_u1299_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({_al_u1794_o,\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o }));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("~(~D*~((C*B))*~(A)+~D*(C*B)*~(A)+~(~D)*(C*B)*A+~D*(C*B)*A)"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0111111100101010),
    .MODE("LOGIC"))
    \_al_u1796|_al_u7150  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [1]}),
    .f({_al_u1796_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0how6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~D)"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b1111111100001111),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u1797|_al_u362  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,open_n9219}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({_al_u1797_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u1800|_al_u909  (
    .b({_al_u909_o,open_n9242}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u1799_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ,_al_u909_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1802|_al_u1648  (
    .a({open_n9263,_al_u1635_o}),
    .b({open_n9264,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u1635_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u1643_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({_al_u1802_o,_al_u1648_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1806|_al_u3792  (
    .a({open_n9289,_al_u1269_o}),
    .b({open_n9290,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u1806_o,_al_u3792_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("(~A*~(D*C*B))"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1808|_al_u1804  (
    .a({_al_u1804_o,_al_u1803_o}),
    .b({_al_u1806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u1808_o,_al_u1804_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1809|_al_u1786  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,open_n9341}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u1296_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u1809_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~(D*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0001000000110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1810|_al_u1811  (
    .a({open_n9362,_al_u1801_o}),
    .b({open_n9363,_al_u1802_o}),
    .c({_al_u1809_o,_al_u1810_o}),
    .d({_al_u1808_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({_al_u1810_o,_al_u1811_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~(~D*~A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*B*~(~D*~A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110000001000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110000001000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1812|_al_u6267  (
    .a({open_n9384,_al_u1385_o}),
    .b({open_n9385,\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u1385_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 }),
    .f({_al_u1812_o,_al_u6267_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1814|_al_u1813  (
    .b({_al_u1813_o,open_n9412}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ,_al_u1813_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1815|_al_u3098  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({_al_u1812_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv }),
    .f({_al_u1815_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u1816|_al_u1582  (
    .b({_al_u1582_o,open_n9467}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u903_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u1816_o,_al_u1582_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1818|_al_u1817  (
    .c({_al_u1817_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u1818_o,_al_u1817_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1819|_al_u605  (
    .a({_al_u1816_o,open_n9516}),
    .b({_al_u1818_o,open_n9517}),
    .c({_al_u604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ,_al_u604_o}),
    .f({_al_u1819_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*C*B*A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000010000000),
    .MODE("LOGIC"))
    \_al_u1820|_al_u1807  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ,open_n9542}),
    .b({_al_u1658_o,open_n9543}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u1820_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(~D*C))"),
    //.LUTF1("(~C*~(B*D))"),
    //.LUTG0("(B*~A*~(~D*C))"),
    //.LUTG1("(~C*~(B*D))"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b0100010000000100),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1822|_al_u1821  (
    .a({open_n9564,_al_u1815_o}),
    .b({_al_u1821_o,_al_u1819_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u1820_o}),
    .d({_al_u1811_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy9iu6 ,_al_u1821_o}));
  // ../RTL/cortexm0ds_logic.v(19971)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1824|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,open_n9589}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ,_al_u1721_o}),
    .f({_al_u1824_o,open_n9604}),
    .q({open_n9608,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 }));  // ../RTL/cortexm0ds_logic.v(19971)
  // ../RTL/cortexm0ds_logic.v(19928)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1827|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,open_n9609}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ,_al_u5103_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 ,_al_u5702_o}),
    .f({_al_u1827_o,open_n9624}),
    .q({open_n9628,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 }));  // ../RTL/cortexm0ds_logic.v(19928)
  // ../RTL/cortexm0ds_logic.v(18358)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1830|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,open_n9629}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cl1iu6 ,open_n9630}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 ,_al_u1753_o}),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ,_al_u1751_o}),
    .f({_al_u1830_o,open_n9645}),
    .q({open_n9649,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 }));  // ../RTL/cortexm0ds_logic.v(18358)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u1832|_al_u4563  (
    .a({\u_cmsdk_mcu/sram_hrdata [17],\u_cmsdk_mcu/sram_hrdata [1]}),
    .b({\u_cmsdk_mcu/flash_hrdata [17],\u_cmsdk_mcu/flash_hrdata [1]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({_al_u1832_o,_al_u4563_o}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1833|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b17  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n9670}),
    .b({_al_u1832_o,open_n9671}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [17]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [17],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1833_o,open_n9684}),
    .q({open_n9688,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [17]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1836|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b18  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n9689}),
    .b({_al_u1835_o,open_n9690}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [18]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1836_o,open_n9707}),
    .q({open_n9711,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [18]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1839|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b19  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n9712}),
    .b({_al_u1838_o,open_n9713}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [19]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [19],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1839_o,open_n9730}),
    .q({open_n9734,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [19]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(B*~(~D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1100110001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1844|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1],open_n9735}),
    .b({_al_u1843_o,_al_u4423_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0],_al_u4438_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u1844_o,\u_cmsdk_mcu/HADDR [2]}),
    .q({open_n9752,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  // ../RTL/cortexm0ds_logic.v(20075)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1846|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6_reg  (
    .a({\u_cmsdk_mcu/sram_hrdata [22],open_n9753}),
    .b({\u_cmsdk_mcu/flash_hrdata [22],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/flash_hrdata [22]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/HWDATA [22]}),
    .mi({open_n9757,\u_cmsdk_mcu/HWDATA [22]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1846_o,\u_cmsdk_mcu/u_ahb_rom/n13 [22]}),
    .q({open_n9772,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 }));  // ../RTL/cortexm0ds_logic.v(20075)
  // ../RTL/cortexm0ds_logic.v(19089)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1848|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6_reg  (
    .a({\u_cmsdk_mcu/sram_hrdata [23],open_n9773}),
    .b({\u_cmsdk_mcu/flash_hrdata [23],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/flash_hrdata [23]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/HWDATA [23]}),
    .mi({open_n9777,\u_cmsdk_mcu/HWDATA [23]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1848_o,\u_cmsdk_mcu/u_ahb_rom/n13 [23]}),
    .q({open_n9792,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 }));  // ../RTL/cortexm0ds_logic.v(19089)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(A*~(~D*C)))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0100010011000100),
    .MODE("LOGIC"))
    \_al_u1859|_al_u1858  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1],\u_cmsdk_mcu/sram_hrdata [28]}),
    .b({_al_u1858_o,\u_cmsdk_mcu/flash_hrdata [28]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({_al_u1859_o,_al_u1858_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1862|_al_u1861  (
    .a({open_n9813,\u_cmsdk_mcu/sram_hrdata [29]}),
    .b({open_n9814,\u_cmsdk_mcu/flash_hrdata [29]}),
    .c({_al_u1861_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({_al_u1862_o,_al_u1861_o}));
  // ../RTL/cortexm0ds_logic.v(19101)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1864|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6_reg  (
    .a({\u_cmsdk_mcu/sram_hrdata [31],open_n9839}),
    .b({\u_cmsdk_mcu/flash_hrdata [31],\u_cmsdk_mcu/sram_hrdata [31]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/HWDATA [31]}),
    .mi({open_n9843,\u_cmsdk_mcu/HWDATA [31]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1864_o,\u_cmsdk_mcu/u_ahb_ram/n13 [31]}),
    .q({open_n9858,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 }));  // ../RTL/cortexm0ds_logic.v(19101)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1868|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b16  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n9859}),
    .b({_al_u1867_o,open_n9860}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [16]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1868_o,open_n9873}),
    .q({open_n9877,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [16]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*~B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"))
    \_al_u1871|_al_u1876  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }));
  // ../RTL/cortexm0ds_logic.v(20177)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1877|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rribx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ,_al_u2414_o}),
    .mi({open_n9905,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ,_al_u2415_o}),
    .q({open_n9921,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[28] }));  // ../RTL/cortexm0ds_logic.v(20177)
  // ../RTL/cortexm0ds_logic.v(18743)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1882|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmlax6_reg  (
    .a({_al_u1875_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N30iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qy2pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1881_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[0] }),
    .mi({open_n9932,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({_al_u1882_o,_al_u1881_o}),
    .q({open_n9937,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] }));  // ../RTL/cortexm0ds_logic.v(18743)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*D))"),
    //.LUT1("(~C*B*~D)"),
    .INIT_LUT0(16'b0000001100001111),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"))
    \_al_u1883|_al_u1892  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .d({_al_u1882_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv }),
    .f({_al_u1883_o,_al_u1892_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1886|_al_u1885  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({_al_u1296_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u1885_o,_al_u914_o}),
    .f({_al_u1886_o,_al_u1885_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1887|_al_u1658  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u1658_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u1887_o,_al_u1658_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1889|_al_u678  (
    .b({_al_u678_o,open_n10012}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ,_al_u678_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1890|_al_u1888  (
    .b({open_n10039,_al_u1887_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u1888_o,_al_u1886_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,_al_u1888_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1891|_al_u2099  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv }),
    .d({_al_u1883_o,_al_u1944_o}),
    .f({_al_u1891_o,_al_u2099_o}));
  // ../RTL/cortexm0ds_logic.v(18867)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1894|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngsax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ,open_n10086}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1893_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv }),
    .mi({open_n10097,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({_al_u1894_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 }),
    .q({open_n10102,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[8] }));  // ../RTL/cortexm0ds_logic.v(18867)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~B*A)"),
    //.LUTF1("(D*~C*~B*A)"),
    //.LUTG0("(D*C*~B*A)"),
    //.LUTG1("(D*~C*~B*A)"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000001000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1897|_al_u1898  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }));
  // ../RTL/cortexm0ds_logic.v(18791)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1900|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9oax6_reg  (
    .a({_al_u1894_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({_al_u1895_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({_al_u1896_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1899_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] }),
    .mi({open_n10130,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({_al_u1900_o,_al_u1896_o}),
    .q({open_n10146,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] }));  // ../RTL/cortexm0ds_logic.v(18791)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1901|_al_u1195  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvzhu6 }),
    .d({_al_u1900_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [8]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~(~D*~A)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100000011000100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1904|_al_u4308  (
    .a({open_n10175,_al_u1643_o}),
    .b({open_n10176,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,_al_u604_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ,_al_u4308_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~B*~(~D*C*A))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~B*~(~D*C*A))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0011001100010011),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0011001100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1906|_al_u1905  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ,open_n10197}),
    .b({_al_u1905_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .c({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 }),
    .f({_al_u1906_o,_al_u1905_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(~D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(~C*B)*~(~D*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111001101010001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001101010001),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1908|_al_u2644  (
    .a({open_n10222,_al_u682_o}),
    .b({open_n10223,_al_u1907_o}),
    .c({_al_u1907_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({_al_u681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv ,_al_u2644_o}));
  // ../RTL/cortexm0ds_logic.v(18848)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1915|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Serax6_reg  (
    .a({_al_u1911_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({_al_u1912_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({_al_u1913_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro2pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 }),
    .mi({open_n10251,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u1915_o,_al_u1912_o}),
    .q({open_n10267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] }));  // ../RTL/cortexm0ds_logic.v(18848)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1916|_al_u5991  (
    .a({open_n10268,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 }),
    .b({open_n10269,_al_u607_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxzhu6 ,_al_u932_o}),
    .d({_al_u1915_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }),
    .f({_al_u1916_o,_al_u5991_o}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1917|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b2  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({_al_u1916_o,_al_u1917_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1917_o,\u_cmsdk_mcu/HWDATA [2]}),
    .q({open_n10311,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [2]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cortexm0ds_logic.v(18744)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1924|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bolax6_reg  (
    .a({_al_u1920_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({_al_u1921_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X62pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1923_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[3] }),
    .mi({open_n10315,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1924_o,_al_u1923_o}),
    .q({open_n10331,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] }));  // ../RTL/cortexm0ds_logic.v(18744)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1925|_al_u1081  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 }),
    .d({_al_u1924_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [3]}));
  // ../RTL/cortexm0ds_logic.v(20152)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1926|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1925_o,_al_u1926_o}),
    .f({_al_u1926_o,\u_cmsdk_mcu/HWDATA [3]}),
    .q({open_n10378,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 }));  // ../RTL/cortexm0ds_logic.v(20152)
  // ../RTL/cortexm0ds_logic.v(18739)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1933|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Delax6_reg  (
    .a({_al_u1929_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({_al_u1930_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kp1pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[4] }),
    .mi({open_n10382,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1933_o,_al_u1930_o}),
    .q({open_n10398,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[4] }));  // ../RTL/cortexm0ds_logic.v(18739)
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*~(D*~B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1000000010100000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1934|_al_u6215  (
    .a({open_n10399,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl4ju6_lutinv }),
    .b({open_n10400,_al_u1934_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwzhu6 ,_al_u6214_o}),
    .d({_al_u1933_o,_al_u5854_o}),
    .f({_al_u1934_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 }));
  // ../RTL/cortexm0ds_logic.v(18875)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1938|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwsax6_reg  (
    .a({open_n10421,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1937_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[5] }),
    .mi({open_n10432,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1938_o,_al_u1937_o}),
    .q({open_n10437,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[5] }));  // ../RTL/cortexm0ds_logic.v(18875)
  // ../RTL/cortexm0ds_logic.v(17288)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1942|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S5kpw6_reg  (
    .a({_al_u1938_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({_al_u1939_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X71pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1941_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] }),
    .mi({open_n10441,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1942_o,_al_u1941_o}),
    .q({open_n10457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[5] }));  // ../RTL/cortexm0ds_logic.v(17288)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1943|_al_u1105  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 }),
    .d({_al_u1942_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1943_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [5]}));
  // ../RTL/cortexm0ds_logic.v(17494)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(~C*B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1944|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1943_o,_al_u1944_o}),
    .f({_al_u1944_o,\u_cmsdk_mcu/HWDATA [5]}),
    .q({open_n10500,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 }));  // ../RTL/cortexm0ds_logic.v(17494)
  // ../RTL/cortexm0ds_logic.v(18746)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1947|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrlax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ,open_n10503}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] ,_al_u5892_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1946_o,_al_u7049_o}),
    .f({_al_u1947_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .q({open_n10520,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[6] }));  // ../RTL/cortexm0ds_logic.v(18746)
  // ../RTL/cortexm0ds_logic.v(18774)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1951|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbnax6_reg  (
    .a({_al_u1947_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({_al_u1948_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq0pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1950_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 }),
    .mi({open_n10531,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1951_o,_al_u1948_o}),
    .q({open_n10536,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[6] }));  // ../RTL/cortexm0ds_logic.v(18774)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1952|_al_u1117  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 }),
    .d({_al_u1951_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1952_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [6]}));
  // ../RTL/cortexm0ds_logic.v(19879)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1953|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1952_o,_al_u1953_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1953_o,\u_cmsdk_mcu/HWDATA [6]}),
    .q({open_n10586,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 }));  // ../RTL/cortexm0ds_logic.v(19879)
  // ../RTL/cortexm0ds_logic.v(18747)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1960|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ytlax6_reg  (
    .a({_al_u1956_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({_al_u1957_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1959_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] }),
    .mi({open_n10597,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u1960_o,_al_u1959_o}),
    .q({open_n10602,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] }));  // ../RTL/cortexm0ds_logic.v(18747)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1961|_al_u1129  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 }),
    .d({_al_u1960_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u1961_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [7]}));
  // ../RTL/cortexm0ds_logic.v(19137)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(~C*B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1962|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1961_o,_al_u1962_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1962_o,\u_cmsdk_mcu/HWDATA [7]}),
    .q({open_n10648,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 }));  // ../RTL/cortexm0ds_logic.v(19137)
  // ../RTL/cortexm0ds_logic.v(18882)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1968|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fatax6_reg  (
    .a({_al_u1965_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O00iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({_al_u1966_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1967_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] }),
    .mi({open_n10659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({_al_u1968_o,_al_u1966_o}),
    .q({open_n10664,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[1] }));  // ../RTL/cortexm0ds_logic.v(18882)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1969|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({_al_u1968_o,_al_u1969_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u1969_o,\u_cmsdk_mcu/HWDATA [1]}),
    .q({open_n10686,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [1]}));  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1971|_al_u2055  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv }),
    .d({_al_u1969_o,_al_u1926_o}),
    .f({_al_u1971_o,_al_u2055_o}));
  // ../RTL/cortexm0ds_logic.v(19772)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1976|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ce7bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] }),
    .mi({open_n10718,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .f({_al_u1976_o,_al_u2056_o}),
    .q({open_n10734,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[11] }));  // ../RTL/cortexm0ds_logic.v(19772)
  // ../RTL/cortexm0ds_logic.v(18866)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1977|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oesax6_reg  (
    .a({_al_u1973_o,open_n10735}),
    .b({_al_u1974_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({_al_u1975_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1976_o,_al_u1972_o}),
    .mi({open_n10746,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({_al_u1977_o,_al_u1973_o}),
    .q({open_n10751,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[9] }));  // ../RTL/cortexm0ds_logic.v(18866)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1978|_al_u1207  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evzhu6 }),
    .d({_al_u1977_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [9]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1981|_al_u1993  (
    .a({open_n10776,_al_u581_o}),
    .b({open_n10777,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6:5]),
    .d({_al_u581_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,_al_u1993_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1982|_al_u1986  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .f({_al_u1982_o,_al_u1986_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u1989|_al_u1988  (
    .b({_al_u588_o,open_n10828}),
    .c({_al_u1988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u1987_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 ,_al_u1988_o}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1991|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b7  (
    .a({_al_u1987_o,open_n10849}),
    .b({_al_u588_o,open_n10850}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n158 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 ,open_n10867}),
    .q({open_n10871,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [7]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1994|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b6  (
    .b({_al_u588_o,open_n10874}),
    .c({_al_u1988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n111 ),
    .clk(XTAL1_wire),
    .d({_al_u1993_o,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 ,open_n10891}),
    .q({open_n10895,\u_cmsdk_mcu/p1_altfunc [6]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1996|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b3  (
    .a({_al_u1993_o,open_n10896}),
    .b({_al_u588_o,open_n10897}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n60 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 ,open_n10910}),
    .q({open_n10914,\u_cmsdk_mcu/p1_outen [3]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2000|_al_u1987  (
    .b({_al_u593_o,open_n10917}),
    .c({_al_u1988_o,_al_u1986_o}),
    .d({_al_u1987_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 ,_al_u1987_o}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2002|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b6  (
    .a({_al_u1987_o,open_n10938}),
    .b({_al_u593_o,open_n10939}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n156 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 ,open_n10952}),
    .q({open_n10956,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [6]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2004|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b6  (
    .b({_al_u593_o,open_n10959}),
    .c({_al_u1988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n111 ),
    .clk(XTAL1_wire),
    .d({_al_u1993_o,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 ,open_n10972}),
    .q({open_n10976,\u_cmsdk_mcu/p0_altfunc [6]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2008|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b0  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],open_n10979}),
    .c({\u_cmsdk_mcu/flash_hrdata [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n99 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [0],open_n10996}),
    .q({open_n11000,\u_cmsdk_mcu/p1_altfunc [0]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2012|_al_u2498  (
    .b({_al_u585_o,_al_u585_o}),
    .c({_al_u1988_o,_al_u1988_o}),
    .d({_al_u1987_o,_al_u1983_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 }));
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2016|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b14  (
    .b({_al_u585_o,open_n11025}),
    .c({_al_u1988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n127 ),
    .clk(XTAL1_wire),
    .d({_al_u1993_o,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 ,open_n11042}),
    .q({open_n11046,\u_cmsdk_mcu/p1_altfunc [14]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2022|_al_u2516  (
    .b({_al_u591_o,_al_u591_o}),
    .c({_al_u1988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u1987_o,_al_u1987_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 ,_al_u2516_o}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2024|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b14  (
    .a({_al_u1987_o,open_n11073}),
    .b({_al_u591_o,open_n11074}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n172 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 ,open_n11087}),
    .q({open_n11091,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [14]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2026|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b14  (
    .b({_al_u591_o,open_n11094}),
    .c({_al_u1988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n127 ),
    .clk(XTAL1_wire),
    .d({_al_u1993_o,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 ,open_n11107}),
    .q({open_n11111,\u_cmsdk_mcu/p0_altfunc [14]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2030|_al_u2628  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]}),
    .c({\u_cmsdk_mcu/flash_hrdata [8],\u_cmsdk_mcu/flash_hrdata [14]}),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [14]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [8],\u_cmsdk_mcu/u_ahb_rom/n13 [14]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2031|_al_u4826  (
    .a({open_n11138,\u_cmsdk_mcu/sram_hrdata [8]}),
    .b({\u_cmsdk_mcu/sram_hrdata [8],\u_cmsdk_mcu/flash_hrdata [8]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [8],_al_u4826_o}));
  // ../RTL/cortexm0ds_logic.v(18890)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2035|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqtax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ,open_n11163}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,_al_u2122_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .mi({open_n11174,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({_al_u2035_o,_al_u2123_o}),
    .q({open_n11179,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[14] }));  // ../RTL/cortexm0ds_logic.v(18890)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u2038|_al_u2034  (
    .a({_al_u2034_o,open_n11180}),
    .b({_al_u2035_o,_al_u2033_o}),
    .c({_al_u2036_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 }),
    .d({_al_u2037_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .f({_al_u2038_o,_al_u2034_o}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2053|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b2  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],open_n11203}),
    .c({\u_cmsdk_mcu/flash_hrdata [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n148 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [2],open_n11220}),
    .q({open_n11224,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [2]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2054|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b2  (
    .b({\u_cmsdk_mcu/sram_hrdata [2],open_n11227}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n103 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [2],open_n11240}),
    .q({open_n11244,\u_cmsdk_mcu/p0_altfunc [2]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cortexm0ds_logic.v(19800)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2061|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zn8bx6_reg  (
    .a({_al_u2057_o,open_n11245}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hy1pw6 ,_al_u2056_o}),
    .c({_al_u2059_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2060_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .mi({open_n11249,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 }),
    .f({_al_u2061_o,_al_u2057_o}),
    .q({open_n11265,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[11] }));  // ../RTL/cortexm0ds_logic.v(19800)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2062|_al_u1087  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z20iu6 }),
    .d({_al_u2061_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2062_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [11]}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2075|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b3  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],open_n11292}),
    .c({\u_cmsdk_mcu/flash_hrdata [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n150 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [3],open_n11309}),
    .q({open_n11313,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [3]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2076|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b3  (
    .b({\u_cmsdk_mcu/sram_hrdata [3],open_n11316}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n105 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [3],open_n11329}),
    .q({open_n11333,\u_cmsdk_mcu/p0_altfunc [3]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2077|_al_u1935  (
    .b({open_n11336,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .d({_al_u1935_o,_al_u1934_o}),
    .f({_al_u2077_o,_al_u1935_o}));
  // ../RTL/cortexm0ds_logic.v(18762)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*B*~D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2082|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnmax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,open_n11361}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ,_al_u7002_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ,_al_u5933_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] ,_al_u6969_o}),
    .f({_al_u2082_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .q({open_n11382,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[12] }));  // ../RTL/cortexm0ds_logic.v(18762)
  // ../RTL/cortexm0ds_logic.v(18864)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2083|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oasax6_reg  (
    .a({_al_u2079_o,open_n11383}),
    .b({_al_u2080_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({_al_u2081_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2082_o,_al_u2078_o}),
    .mi({open_n11387,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u2083_o,_al_u2079_o}),
    .q({open_n11403,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[12] }));  // ../RTL/cortexm0ds_logic.v(18864)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2084|_al_u1099  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S20iu6 }),
    .d({_al_u2083_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2084_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [12]}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2097|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b4  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],open_n11434}),
    .c({\u_cmsdk_mcu/flash_hrdata [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n152 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [4],open_n11451}),
    .q({open_n11455,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [4]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2098|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b4  (
    .b({\u_cmsdk_mcu/sram_hrdata [4],open_n11458}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n107 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [4],open_n11475}),
    .q({open_n11479,\u_cmsdk_mcu/p1_altfunc [4]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cortexm0ds_logic.v(17301)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2105|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlkpw6_reg  (
    .a({_al_u2101_o,open_n11480}),
    .b({_al_u2102_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2104_o,_al_u2100_o}),
    .mi({open_n11491,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({_al_u2105_o,_al_u2101_o}),
    .q({open_n11496,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] }));  // ../RTL/cortexm0ds_logic.v(17301)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2106|_al_u1111  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L20iu6 }),
    .d({_al_u2105_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2106_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [13]}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2119|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b5  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],open_n11527}),
    .c({\u_cmsdk_mcu/flash_hrdata [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n64 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [5],open_n11540}),
    .q({open_n11544,\u_cmsdk_mcu/p1_outen [5]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b5  (
    .b({\u_cmsdk_mcu/sram_hrdata [5],open_n11547}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n154 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [5],open_n11564}),
    .q({open_n11568,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [5]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cortexm0ds_logic.v(19569)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~A*~(~C*B))"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110101110),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2121|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6_reg  (
    .a({open_n11569,_al_u2121_o}),
    .b({open_n11570,_al_u1892_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,_al_u2128_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1953_o,_al_u2129_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2121_o,\u_cmsdk_mcu/HWDATA [14]}),
    .q({open_n11586,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 }));  // ../RTL/cortexm0ds_logic.v(19569)
  // ../RTL/cortexm0ds_logic.v(18115)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2127|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S38ax6_reg  (
    .a({_al_u2123_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({_al_u2124_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({_al_u2125_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2126_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] }),
    .mi({open_n11590,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({_al_u2127_o,_al_u2125_o}),
    .q({open_n11606,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[14] }));  // ../RTL/cortexm0ds_logic.v(18115)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2128|_al_u1123  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E20iu6 }),
    .d({_al_u2127_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2128_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [14]}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~A*~(~C*B))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110101110),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2143|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b15  (
    .a({open_n11631,_al_u2143_o}),
    .b({open_n11632,_al_u1892_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,_al_u2150_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({_al_u1962_o,_al_u2151_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2143_o,\u_cmsdk_mcu/HWDATA [15]}),
    .q({open_n11648,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [15]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cortexm0ds_logic.v(19789)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2149|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18bx6_reg  (
    .a({_al_u2145_o,open_n11649}),
    .b({_al_u2146_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2148_o,_al_u2144_o}),
    .mi({open_n11653,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u2149_o,_al_u2145_o}),
    .q({open_n11669,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[15] }));  // ../RTL/cortexm0ds_logic.v(19789)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2150|_al_u1135  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X10iu6 }),
    .d({_al_u2149_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2150_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [15]}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2163|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b7  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],open_n11696}),
    .c({\u_cmsdk_mcu/flash_hrdata [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n158 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [7],open_n11709}),
    .q({open_n11713,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [7]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2164|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b7  (
    .b({\u_cmsdk_mcu/sram_hrdata [7],open_n11716}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n113 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [7],open_n11733}),
    .q({open_n11737,\u_cmsdk_mcu/p1_altfunc [7]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cortexm0ds_logic.v(18860)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2170|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2sax6_reg  (
    .a({_al_u2166_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({_al_u2167_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({_al_u2168_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drzow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 }),
    .mi({open_n11741,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u2170_o,_al_u2167_o}),
    .q({open_n11757,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[17] }));  // ../RTL/cortexm0ds_logic.v(18860)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2171|_al_u1141  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J10iu6 }),
    .d({_al_u2170_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2171_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2172|_al_u2174  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .d({_al_u1888_o,_al_u1888_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2187|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b1  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],open_n11814}),
    .c({\u_cmsdk_mcu/flash_hrdata [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n146 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [1],open_n11831}),
    .q({open_n11835,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [1]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2188|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b1  (
    .b({\u_cmsdk_mcu/sram_hrdata [1],open_n11838}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n101 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [1],open_n11851}),
    .q({open_n11855,\u_cmsdk_mcu/p0_altfunc [1]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2199|_al_u2580  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]}),
    .c({\u_cmsdk_mcu/flash_hrdata [9],\u_cmsdk_mcu/flash_hrdata [12]}),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [12]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [9],\u_cmsdk_mcu/u_ahb_rom/n13 [12]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2200|_al_u2663  (
    .b({\u_cmsdk_mcu/sram_hrdata [9],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/flash_hrdata [15]}),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [15]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [9],\u_cmsdk_mcu/u_ahb_rom/n13 [15]}));
  // ../RTL/cortexm0ds_logic.v(18887)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2207|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ektax6_reg  (
    .a({_al_u2203_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({_al_u2204_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({_al_u2205_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eazow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] }),
    .mi({open_n11914,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u2207_o,_al_u2205_o}),
    .q({open_n11919,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[18] }));  // ../RTL/cortexm0ds_logic.v(18887)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2208|_al_u1153  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10iu6 }),
    .d({_al_u2207_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2208_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [18]}));
  // ../RTL/cortexm0ds_logic.v(18756)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2212|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbmax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2211_o,_al_u6844_o}),
    .f({_al_u2212_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .q({open_n11962,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[19] }));  // ../RTL/cortexm0ds_logic.v(18756)
  // ../RTL/cortexm0ds_logic.v(17782)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2216|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jtvpw6_reg  (
    .a({_al_u2212_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgqow6 }),
    .b({_al_u2213_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2215_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] }),
    .mi({open_n11966,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({_al_u2216_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zow6 }),
    .q({open_n11982,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[17] }));  // ../RTL/cortexm0ds_logic.v(17782)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2217|_al_u1159  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V00iu6 }),
    .d({_al_u2216_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2217_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [19]}));
  // ../RTL/cortexm0ds_logic.v(18755)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2224|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9max6_reg  (
    .a({_al_u2220_o,open_n12011}),
    .b({_al_u2221_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqyow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2223_o,_al_u2219_o}),
    .mi({open_n12022,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .f({_al_u2224_o,_al_u2220_o}),
    .q({open_n12027,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[20] }));  // ../RTL/cortexm0ds_logic.v(18755)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2225|_al_u1165  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H00iu6 }),
    .d({_al_u2224_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [20]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u2234|_al_u2230  (
    .a({_al_u2230_o,open_n12056}),
    .b({_al_u2231_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhyow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] }),
    .d({_al_u2233_o,_al_u2229_o}),
    .f({_al_u2234_o,_al_u2230_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2235|_al_u1171  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A00iu6 }),
    .d({_al_u2234_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2235_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [21]}));
  // ../RTL/cortexm0ds_logic.v(20009)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2239|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tbfbx6_reg  (
    .a({open_n12101,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2238_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] }),
    .mi({open_n12105,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u2239_o,_al_u2238_o}),
    .q({open_n12121,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[22] }));  // ../RTL/cortexm0ds_logic.v(20009)
  // ../RTL/cortexm0ds_logic.v(20001)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2243|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tvebx6_reg  (
    .a({_al_u2239_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({_al_u2240_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7yow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2242_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] }),
    .mi({open_n12132,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u2243_o,_al_u2242_o}),
    .q({open_n12137,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] }));  // ../RTL/cortexm0ds_logic.v(20001)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2244|_al_u1177  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzzhu6 }),
    .d({_al_u2243_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2244_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [22]}));
  // ../RTL/cortexm0ds_logic.v(18063)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2251|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P54qw6_reg  (
    .a({_al_u2247_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({_al_u2248_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyxow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2250_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[23] }),
    .mi({open_n12172,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u2251_o,_al_u2250_o}),
    .q({open_n12177,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[23] }));  // ../RTL/cortexm0ds_logic.v(18063)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2252|_al_u1183  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzzhu6 }),
    .d({_al_u2251_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2252_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [23]}));
  // ../RTL/cortexm0ds_logic.v(18855)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2260|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Osrax6_reg  (
    .a({_al_u2256_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({_al_u2257_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6xow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2259_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[25] }),
    .mi({open_n12216,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u2260_o,_al_u2259_o}),
    .q({open_n12221,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[25] }));  // ../RTL/cortexm0ds_logic.v(18855)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2261|_al_u1201  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yyzhu6 }),
    .d({_al_u2260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2261_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [25]}));
  // ../RTL/cortexm0ds_logic.v(17889)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2262|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npypw6_reg  (
    .a({_al_u2261_o,open_n12246}),
    .b({_al_u1968_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] }),
    .c({_al_u1906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkliu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1299_o,_al_u2262_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2262_o,open_n12263}),
    .q({open_n12267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o }));  // ../RTL/cortexm0ds_logic.v(17889)
  // ../RTL/cortexm0ds_logic.v(18769)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2269|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1nax6_reg  (
    .a({_al_u2265_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .b({_al_u2266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .c({_al_u2267_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2268_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] }),
    .mi({open_n12271,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({_al_u2269_o,_al_u2266_o}),
    .q({open_n12287,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[30] }));  // ../RTL/cortexm0ds_logic.v(18769)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2270|_al_u1231  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixzhu6 }),
    .d({_al_u2269_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2270_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [30]}));
  // ../RTL/cortexm0ds_logic.v(18742)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2276|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cklax6_reg  (
    .a({open_n12312,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({_al_u2275_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[31] }),
    .mi({open_n12323,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u2276_o,_al_u2275_o}),
    .q({open_n12328,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[31] }));  // ../RTL/cortexm0ds_logic.v(18742)
  // ../RTL/cortexm0ds_logic.v(18872)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2280|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqsax6_reg  (
    .a({_al_u2276_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({_al_u2277_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({_al_u2278_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2279_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[31] }),
    .mi({open_n12339,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u2280_o,_al_u2278_o}),
    .q({open_n12344,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[31] }));  // ../RTL/cortexm0ds_logic.v(18872)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2281|_al_u1237  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxzhu6 }),
    .d({_al_u2280_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2281_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [31]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2289|_al_u1249  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q10iu6 }),
    .d({_al_u2288_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2289_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~D*~(C@B))"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~D*~(C@B))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000011000011),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000011000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2293|_al_u2292  (
    .a({open_n12393,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .d({_al_u2292_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 }),
    .f({_al_u2293_o,_al_u2292_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~B*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000100000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2295|_al_u2294  (
    .a({open_n12418,_al_u1250_o}),
    .b({open_n12419,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .d({_al_u2293_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .f({_al_u2295_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 }));
  // ../RTL/cortexm0ds_logic.v(17356)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*A)))"),
    //.LUT1("(~A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111100001111),
    .INIT_LUT1(16'b0001010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2297|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6_reg  (
    .a({_al_u2295_o,_al_u2297_o}),
    .b({_al_u2296_o,_al_u2306_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Spyhu6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rsyhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u2297_o,open_n12453}),
    .q({open_n12457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }));  // ../RTL/cortexm0ds_logic.v(17356)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2299|_al_u2298  (
    .b({_al_u2298_o,open_n12460}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .d({_al_u1250_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .f({_al_u2299_o,_al_u2298_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~A*~(D*C*B))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2301|_al_u2300  (
    .a({_al_u2299_o,open_n12485}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ,open_n12486}),
    .c({_al_u1251_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2303|_al_u4027  (
    .b({open_n12513,_al_u3390_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .d({_al_u1757_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ,_al_u4027_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2304|_al_u2302  (
    .b({open_n12540,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 ,_al_u529_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2309|_al_u5211  (
    .b({open_n12567,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azeiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fviow6 }),
    .f({_al_u2309_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yuiow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u2310|_al_u2313  (
    .a({_al_u2309_o,_al_u2309_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozeiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }));
  // ../RTL/cortexm0ds_logic.v(20046)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2315|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n12612}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [22]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ,_al_u2315_o}),
    .f({_al_u2315_o,open_n12631}),
    .q({open_n12635,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 }));  // ../RTL/cortexm0ds_logic.v(20046)
  // ../RTL/cortexm0ds_logic.v(17300)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2317|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12636}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [21],_al_u2317_o}),
    .f({_al_u2317_o,open_n12651}),
    .q({open_n12655,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 }));  // ../RTL/cortexm0ds_logic.v(17300)
  // ../RTL/cortexm0ds_logic.v(17231)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2319|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12656}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [20],_al_u2319_o}),
    .f({_al_u2319_o,open_n12671}),
    .q({open_n12675,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 }));  // ../RTL/cortexm0ds_logic.v(17231)
  // ../RTL/cortexm0ds_logic.v(18109)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2321|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n12676}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [19]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 ,_al_u2321_o}),
    .f({_al_u2321_o,open_n12695}),
    .q({open_n12699,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 }));  // ../RTL/cortexm0ds_logic.v(18109)
  // ../RTL/cortexm0ds_logic.v(17829)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2323|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12700}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [18],_al_u2323_o}),
    .f({_al_u2323_o,open_n12719}),
    .q({open_n12723,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 }));  // ../RTL/cortexm0ds_logic.v(17829)
  // ../RTL/cortexm0ds_logic.v(17710)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2325|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12724}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [17],_al_u2325_o}),
    .f({_al_u2325_o,open_n12739}),
    .q({open_n12743,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 }));  // ../RTL/cortexm0ds_logic.v(17710)
  // ../RTL/cortexm0ds_logic.v(17659)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2327|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12744}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [16],_al_u2327_o}),
    .f({_al_u2327_o,open_n12759}),
    .q({open_n12763,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 }));  // ../RTL/cortexm0ds_logic.v(17659)
  // ../RTL/cortexm0ds_logic.v(18960)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2329|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12764}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [15],_al_u2329_o}),
    .f({_al_u2329_o,open_n12779}),
    .q({open_n12783,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 }));  // ../RTL/cortexm0ds_logic.v(18960)
  // ../RTL/cortexm0ds_logic.v(18961)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2331|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n12784}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,open_n12785}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 ,_al_u2512_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({open_n12789,\u_cmsdk_mcu/HWDATA [14]}),
    .f({_al_u2331_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n262 }),
    .q({open_n12805,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 }));  // ../RTL/cortexm0ds_logic.v(18961)
  // ../RTL/cortexm0ds_logic.v(17290)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2333|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12806}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [13],_al_u2333_o}),
    .f({_al_u2333_o,open_n12821}),
    .q({open_n12825,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 }));  // ../RTL/cortexm0ds_logic.v(17290)
  // ../RTL/cortexm0ds_logic.v(17227)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2335|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12826}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [12],_al_u2335_o}),
    .f({_al_u2335_o,open_n12845}),
    .q({open_n12849,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 }));  // ../RTL/cortexm0ds_logic.v(17227)
  // ../RTL/cortexm0ds_logic.v(18110)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2337|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12850}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [11],_al_u2337_o}),
    .f({_al_u2337_o,open_n12869}),
    .q({open_n12873,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 }));  // ../RTL/cortexm0ds_logic.v(18110)
  // ../RTL/cortexm0ds_logic.v(17689)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~A*~(~C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~D*~A*~(~C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110101110),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111111110101110),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2339|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,_al_u2032_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,_al_u1892_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ,_al_u2040_o}),
    .f({_al_u2339_o,\u_cmsdk_mcu/HWDATA [10]}),
    .q({open_n12894,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 }));  // ../RTL/cortexm0ds_logic.v(17689)
  // ../RTL/cortexm0ds_logic.v(20209)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2341|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12895}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [9],_al_u2341_o}),
    .f({_al_u2341_o,open_n12914}),
    .q({open_n12918,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 }));  // ../RTL/cortexm0ds_logic.v(20209)
  // ../RTL/cortexm0ds_logic.v(17927)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~A*~(~C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~D*~A*~(~C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110101110),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111111110101110),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2343|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,_al_u1891_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,_al_u1892_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 ,_al_u1902_o}),
    .f({_al_u2343_o,\u_cmsdk_mcu/HWDATA [8]}),
    .q({open_n12939,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 }));  // ../RTL/cortexm0ds_logic.v(17927)
  // ../RTL/cortexm0ds_logic.v(18963)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2345|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n12940}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,open_n12941}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 ,_al_u2478_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n12945,\u_cmsdk_mcu/HWDATA [7]}),
    .f({_al_u2345_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n203 }),
    .q({open_n12961,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 }));  // ../RTL/cortexm0ds_logic.v(18963)
  // ../RTL/cortexm0ds_logic.v(18111)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2347|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n12962}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [6],_al_u2347_o}),
    .f({_al_u2347_o,open_n12981}),
    .q({open_n12985,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 }));  // ../RTL/cortexm0ds_logic.v(18111)
  // ../RTL/cortexm0ds_logic.v(17495)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2349|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n12986}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [5]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ,_al_u2349_o}),
    .f({_al_u2349_o,open_n13005}),
    .q({open_n13009,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 }));  // ../RTL/cortexm0ds_logic.v(17495)
  // ../RTL/cortexm0ds_logic.v(20127)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2351|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n13010}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [4],_al_u2351_o}),
    .f({_al_u2351_o,open_n13025}),
    .q({open_n13029,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 }));  // ../RTL/cortexm0ds_logic.v(20127)
  // ../RTL/cortexm0ds_logic.v(20153)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2353|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n13030}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [3]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ,_al_u2353_o}),
    .f({_al_u2353_o,open_n13045}),
    .q({open_n13049,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 }));  // ../RTL/cortexm0ds_logic.v(20153)
  // ../RTL/cortexm0ds_logic.v(19903)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2355|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,open_n13050}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [2],_al_u2355_o}),
    .f({_al_u2355_o,open_n13069}),
    .q({open_n13073,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 }));  // ../RTL/cortexm0ds_logic.v(19903)
  // ../RTL/cortexm0ds_logic.v(18966)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2357|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n13074}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,open_n13075}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 ,\u_cmsdk_mcu/HWDATA [1]}),
    .f({_al_u2357_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 }),
    .q({open_n13092,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 }));  // ../RTL/cortexm0ds_logic.v(18966)
  // ../RTL/cortexm0ds_logic.v(17599)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2359|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv ,open_n13093}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [0]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 ,_al_u2359_o}),
    .f({_al_u2359_o,open_n13108}),
    .q({open_n13112,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 }));  // ../RTL/cortexm0ds_logic.v(17599)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2362|_al_u911  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ,open_n13115}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u2361_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u2363|_al_u2767  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({_al_u1812_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,_al_u2767_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2365|_al_u2364  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u2364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({_al_u2365_o,_al_u2364_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2366|_al_u4037  (
    .a({_al_u1802_o,open_n13192}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 ,_al_u3227_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u2365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv }),
    .f({_al_u2366_o,_al_u4037_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2368|_al_u2367  (
    .c({_al_u2367_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ,_al_u2367_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*A*~(~D*B))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(~C*A*~(~D*B))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0000101000000010),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2372|_al_u2370  (
    .a({_al_u2366_o,_al_u2369_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({_al_u2370_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u2371_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ,_al_u2370_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2374|_al_u2373  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,open_n13271}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u2373_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhow6 ,_al_u2373_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2376|_al_u1369  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u2376_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~D*~C*B))"),
    //.LUT1("(~B*A*~(~D*C))"),
    .INIT_LUT0(16'b0101010101010001),
    .INIT_LUT1(16'b0010001000000010),
    .MODE("LOGIC"))
    \_al_u2377|_al_u2375  (
    .a({_al_u2375_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhow6 }),
    .b({_al_u2376_o,_al_u2364_o}),
    .c({_al_u2364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u2377_o,_al_u2375_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(A*~(D*~C*~B))"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(A*~(D*~C*~B))"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b1010100010101010),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b1010100010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2379|_al_u2378  (
    .a({_al_u2377_o,open_n13340}),
    .b({_al_u2378_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({_al_u2379_o,_al_u2378_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2382|_al_u2381  (
    .a({_al_u2379_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 }),
    .b({_al_u1815_o,_al_u2380_o}),
    .c({_al_u2361_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({_al_u2381_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({_al_u2382_o,_al_u2381_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2385|_al_u2384  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~(~D*A)))"),
    //.LUTF1("(~C*~(B*D))"),
    //.LUTG0("(C*~(~B*~(~D*A)))"),
    //.LUTG1("(~C*~(B*D))"),
    .INIT_LUTF0(16'b1100000011100000),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b1100000011100000),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2389|_al_u2388  (
    .a({open_n13413,_al_u932_o}),
    .b({_al_u2386_o,_al_u2387_o}),
    .c({_al_u2388_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u2389_o,_al_u2388_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~D*~C*A))"),
    //.LUTF1("~(~D*~(C*B*A))"),
    //.LUTG0("(B*~(~D*~C*A))"),
    //.LUTG1("~(~D*~(C*B*A))"),
    .INIT_LUTF0(16'b1100110011000100),
    .INIT_LUTF1(16'b1111111110000000),
    .INIT_LUTG0(16'b1100110011000100),
    .INIT_LUTG1(16'b1111111110000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2391|_al_u2390  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 }),
    .b({_al_u2382_o,_al_u2389_o}),
    .c({_al_u2390_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ,_al_u2390_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(~D*C))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(B*A*~(~D*C))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1000100000001000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1000100000001000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2393|_al_u3819  (
    .a({open_n13462,_al_u903_o}),
    .b({_al_u1583_o,_al_u2392_o}),
    .c({_al_u2392_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u1663_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .f({_al_u2393_o,_al_u3819_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(D*(C@B))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0011110000000000),
    .MODE("LOGIC"))
    \_al_u2395|_al_u2394  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,open_n13489}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u2395_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2396|_al_u1662  (
    .b({_al_u1662_o,open_n13512}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u2396_o,_al_u1662_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b1011111110110011),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1011111110110011),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2397|_al_u2440  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lu0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 }),
    .b({_al_u2393_o,_al_u2413_o}),
    .c({_al_u2395_o,_al_u2439_o}),
    .d({_al_u2396_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv }),
    .f({_al_u2397_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUT1("(C*~(~B*~D))"),
    .INIT_LUT0(16'b0001111100110101),
    .INIT_LUT1(16'b1111000011000000),
    .MODE("LOGIC"))
    \_al_u2401|_al_u3008  (
    .a({open_n13561,_al_u2399_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 }),
    .d({_al_u2399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv ,_al_u3008_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D)*~(B)*~(C)+~(D)*B*~(C)+D*B*~(C)+D*~(B)*C+D*B*C)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111110000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2402|_al_u2413  (
    .b({open_n13584,_al_u2412_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk8ju6_lutinv }),
    .d({_al_u2398_o,_al_u2398_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,_al_u2413_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2404|_al_u2403  (
    .b({_al_u2403_o,open_n13607}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u2404_o,_al_u2403_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2407|_al_u2406  (
    .b({_al_u2406_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u695_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u2407_o,_al_u2406_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~A*~(~D*~(~C*~B)))"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0101010100000001),
    .MODE("LOGIC"))
    \_al_u2411|_al_u2409  (
    .a({_al_u2409_o,open_n13658}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv }),
    .f({_al_u2411_o,_al_u2409_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(C*B)))"),
    //.LUT1("(D*~(C*~B*~A))"),
    .INIT_LUT0(16'b1110101000000000),
    .INIT_LUT1(16'b1110111100000000),
    .MODE("LOGIC"))
    \_al_u2412|_al_u2405  (
    .a({_al_u2405_o,_al_u2404_o}),
    .b({_al_u2407_o,_al_u604_o}),
    .c({_al_u2411_o,_al_u1344_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u2412_o,_al_u2405_o}));
  // ../RTL/cortexm0ds_logic.v(20169)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2419|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rbibx6_reg  (
    .a({_al_u2415_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({_al_u2416_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({_al_u2417_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2418_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[28] }),
    .mi({open_n13709,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({_al_u2419_o,_al_u2418_o}),
    .q({open_n13714,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[28] }));  // ../RTL/cortexm0ds_logic.v(20169)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2420|_al_u1225  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyzhu6 }),
    .d({_al_u2419_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2420_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [28]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2421|_al_u2398  (
    .c({_al_u2412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .d({_al_u2397_o,_al_u2397_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,_al_u2398_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1011111110110011),
    .MODE("LOGIC"))
    \_al_u2422|_al_u1526  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,open_n13771}),
    .b({_al_u2413_o,open_n13772}),
    .c({_al_u2420_o,_al_u1348_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,_al_u1525_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [28]}));
  // ../RTL/cortexm0ds_logic.v(17247)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2428|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkjpw6_reg  (
    .a({_al_u2424_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({_al_u2425_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({_al_u2426_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2427_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] }),
    .mi({open_n13803,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u2428_o,_al_u2426_o}),
    .q({open_n13808,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[29] }));  // ../RTL/cortexm0ds_logic.v(17247)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2429|_al_u1243  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxzhu6 }),
    .d({_al_u2428_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2429_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [29]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(~B*A))"),
    //.LUTF1("~(B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUTG0("(~(D*C)*~(~B*A))"),
    //.LUTG1("~(B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT_LUTF0(16'b0000110111011101),
    .INIT_LUTF1(16'b1011101111110011),
    .INIT_LUTG0(16'b0000110111011101),
    .INIT_LUTG1(16'b1011101111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2430|_al_u2740  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .b({_al_u2413_o,_al_u2429_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 }),
    .d({_al_u2429_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29],_al_u2740_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("~(C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("~(C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b1101111110001111),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b1101111110001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2431|_al_u5859  (
    .a({_al_u2270_o,open_n13861}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,_al_u5858_o}),
    .c({_al_u2413_o,_al_u5854_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,_al_u2270_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30],_al_u5859_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*C*A))"),
    //.LUTF1("~(C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    //.LUTG0("(B*~(D*C*A))"),
    //.LUTG1("~(C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT_LUTF0(16'b0100110011001100),
    .INIT_LUTF1(16'b1101111110001111),
    .INIT_LUTG0(16'b0100110011001100),
    .INIT_LUTG1(16'b1101111110001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2432|_al_u5870  (
    .a({_al_u2261_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,_al_u5869_o}),
    .c({_al_u2413_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25],_al_u5870_o}));
  // ../RTL/cortexm0ds_logic.v(18776)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2438|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfnax6_reg  (
    .a({_al_u2434_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({_al_u2435_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voxow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2437_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[24] }),
    .mi({open_n13913,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u2438_o,_al_u2435_o}),
    .q({open_n13929,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[24] }));  // ../RTL/cortexm0ds_logic.v(18776)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2439|_al_u1189  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzzhu6 }),
    .d({_al_u2438_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2439_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [24]}));
  // ../RTL/cortexm0ds_logic.v(18778)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2446|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njnax6_reg  (
    .a({_al_u2442_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({_al_u2443_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdwow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2445_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[27] }),
    .mi({open_n13968,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u2446_o,_al_u2443_o}),
    .q({open_n13973,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] }));  // ../RTL/cortexm0ds_logic.v(18778)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2447|_al_u1219  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kyzhu6 }),
    .d({_al_u2446_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2447_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [27]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*C*A))"),
    //.LUT1("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT_LUT0(16'b0100110011001100),
    .INIT_LUT1(16'b1011111110110011),
    .MODE("LOGIC"))
    \_al_u2448|_al_u5905  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27]}),
    .b({_al_u2413_o,_al_u5904_o}),
    .c({_al_u2447_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27],_al_u5905_o}));
  // ../RTL/cortexm0ds_logic.v(17696)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2454|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X3upw6_reg  (
    .a({_al_u2450_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .b({_al_u2451_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynwow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2453_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[26] }),
    .mi({open_n14032,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u2454_o,_al_u2453_o}),
    .q({open_n14037,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[26] }));  // ../RTL/cortexm0ds_logic.v(17696)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2455|_al_u1213  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryzhu6 }),
    .d({_al_u2454_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u2455_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [26]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*C*A))"),
    //.LUTF1("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG0("(B*~(D*C*A))"),
    //.LUTG1("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT_LUTF0(16'b0100110011001100),
    .INIT_LUTF1(16'b1011111110110011),
    .INIT_LUTG0(16'b0100110011001100),
    .INIT_LUTG1(16'b1011111110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2456|_al_u5910  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26]}),
    .b({_al_u2413_o,_al_u5909_o}),
    .c({_al_u2455_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26],_al_u5910_o}));
  // ../RTL/cortexm0ds_logic.v(19029)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~A*~(~D*C))"),
    //.LUT1("~(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101111111011),
    .INIT_LUT1(16'b1011111110110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2457|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T75ju6 ,_al_u2143_o}),
    .b({_al_u2413_o,_al_u2274_o}),
    .c({_al_u2281_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A85ju6_lutinv ,_al_u2281_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ,\u_cmsdk_mcu/HWDATA [31]}),
    .q({open_n14101,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 }));  // ../RTL/cortexm0ds_logic.v(19029)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*B*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"))
    \_al_u2458|_al_u699  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,open_n14104}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u2458_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(A*~(~D*C*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(A*~(~D*C*B))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1010101000101010),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1010101000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2460|_al_u1342  (
    .a({_al_u2459_o,open_n14125}),
    .b({_al_u1342_o,open_n14126}),
    .c({_al_u2403_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u2460_o,_al_u1342_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*A*~(D*C))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*A*~(D*C))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000001000100010),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2462|_al_u2461  (
    .a({open_n14151,_al_u2460_o}),
    .b({open_n14152,_al_u1820_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .d({_al_u2461_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ,_al_u2461_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u2464|_al_u2463  (
    .a({open_n14177,_al_u2399_o}),
    .b({_al_u2463_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({_al_u2464_o,_al_u2463_o}));
  // ../RTL/cortexm0ds_logic.v(17180)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2466|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf1iu6 }),
    .q({open_n14218,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3ipw6 }));  // ../RTL/cortexm0ds_logic.v(17180)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u2467|_al_u3774  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 ,open_n14219}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ,open_n14220}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 }),
    .f({_al_u2467_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*~(C*B)))"),
    //.LUT1("(~D*B*~(C*A))"),
    .INIT_LUT0(16'b1010101010000000),
    .INIT_LUT1(16'b0000000001001100),
    .MODE("LOGIC"))
    \_al_u2469|_al_u1672  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gf1ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 }),
    .f({_al_u2469_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2472|_al_u1048  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ,open_n14263}),
    .c({_al_u1048_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .d({_al_u473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ,_al_u1048_o}));
  // ../RTL/cmsdk_apb_uart.v(634)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("~(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b1111110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2473|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_txintr_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [0],uart0_txen_pad}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n114 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],_al_u637_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n114 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [0]}),
    .q({open_n14301,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]}));  // ../RTL/cmsdk_apb_uart.v(634)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2474|_al_u1983  (
    .b({_al_u588_o,open_n14304}),
    .c({_al_u1988_o,_al_u1982_o}),
    .d({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,_al_u1983_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2475|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b0  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,open_n14331}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n271 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n271 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [0]}),
    .q({open_n14347,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2476|_al_u1984  (
    .a({open_n14348,_al_u1983_o}),
    .b({_al_u588_o,_al_u588_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }));
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2477|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b0  (
    .c({_al_u2476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n234 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n234 ,open_n14393}),
    .q({open_n14397,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [0]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2478|_al_u2480  (
    .b({_al_u588_o,_al_u588_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u1987_o,_al_u1987_o}),
    .f({_al_u2478_o,_al_u2480_o}));
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2479|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b0  (
    .c({_al_u2478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n189 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n189 ,open_n14444}),
    .q({open_n14448,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2481|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b0  (
    .c({_al_u2480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n144 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n144 ,open_n14465}),
    .q({open_n14469,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [0]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2482|_al_u2484  (
    .b({_al_u588_o,_al_u588_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u1993_o,_al_u1993_o}),
    .f({_al_u2482_o,_al_u2484_o}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2483|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b5  (
    .c({_al_u2482_o,_al_u2482_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [5]}),
    .mi({open_n14506,\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n99 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n109 }),
    .q({open_n14510,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [5]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2485|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b6  (
    .c({_al_u2484_o,_al_u2484_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n14525,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n54 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n66 }),
    .q({open_n14529,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [6]}));  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2486|_al_u2510  (
    .b({_al_u593_o,_al_u591_o}),
    .c({_al_u1988_o,_al_u1988_o}),
    .d({_al_u1983_o,_al_u1983_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 }));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2487|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b0  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n271 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n271 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [0]}),
    .q({open_n14573,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2488|_al_u1998  (
    .a({open_n14574,_al_u1983_o}),
    .b({_al_u593_o,_al_u593_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2488_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }));
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2489|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b0  (
    .c({_al_u2488_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n234 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n234 ,open_n14619}),
    .q({open_n14623,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [0]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2490|_al_u2496  (
    .b({_al_u593_o,_al_u593_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u1987_o,_al_u1993_o}),
    .f({_al_u2490_o,_al_u2496_o}));
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2491|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b0  (
    .c({_al_u2490_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n189 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n189 ,open_n14666}),
    .q({open_n14670,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [0]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2492|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b4  (
    .b({_al_u593_o,open_n14673}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4]}),
    .clk(1'b1),
    .d({_al_u1987_o,_al_u3058_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2492_o,open_n14691}),
    .q({open_n14695,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [4]}));  // ../RTL/gpio_ctrl.v(248)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2493|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b0  (
    .c({_al_u2492_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n144 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n144 ,open_n14712}),
    .q({open_n14716,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [0]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2494|_al_u2006  (
    .a({open_n14717,_al_u1993_o}),
    .b({_al_u593_o,_al_u593_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1993_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2494_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }));
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2495|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b0  (
    .c({_al_u2494_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n99 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n99 ,open_n14758}),
    .q({open_n14762,\u_cmsdk_mcu/p0_altfunc [0]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2497|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b0  (
    .c({_al_u2496_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n54 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n54 ,open_n14779}),
    .q({open_n14783,\u_cmsdk_mcu/p0_outen [0]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2499|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b8  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n14786}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n287 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n287 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [8]}),
    .q({open_n14806,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u2500|_al_u2010  (
    .a({open_n14807,_al_u1983_o}),
    .b({_al_u585_o,_al_u585_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }));
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2501|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b8  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n250 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n250 ,open_n14848}),
    .q({open_n14852,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [8]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2502|_al_u2014  (
    .a({open_n14853,_al_u1987_o}),
    .b({_al_u585_o,_al_u585_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1987_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }));
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2503|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b8  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n205 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n205 ,open_n14898}),
    .q({open_n14902,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2504|_al_u2508  (
    .b({_al_u585_o,_al_u585_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u1987_o,_al_u1993_o}),
    .f({_al_u2504_o,_al_u2508_o}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2505|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b8  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n160 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n160 ,open_n14945}),
    .q({open_n14949,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [8]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2506|_al_u2018  (
    .a({open_n14950,_al_u1993_o}),
    .b({_al_u585_o,_al_u585_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1993_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }));
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2507|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b8  (
    .c({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n115 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n115 ,open_n14991}),
    .q({open_n14995,\u_cmsdk_mcu/p1_altfunc [8]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2509|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b8  (
    .c({_al_u2508_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n70 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n70 ,open_n15012}),
    .q({open_n15016,\u_cmsdk_mcu/p1_outen [8]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2511|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b8  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [8]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n287 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n287 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [8]}),
    .q({open_n15034,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u2512|_al_u2020  (
    .a({open_n15035,_al_u1983_o}),
    .b({_al_u591_o,_al_u591_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }));
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2513|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b8  (
    .c({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n250 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n250 ,open_n15076}),
    .q({open_n15080,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [8]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2514|_al_u2520  (
    .b({_al_u591_o,_al_u591_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u1987_o,_al_u1993_o}),
    .f({_al_u2514_o,_al_u2520_o}));
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2515|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b8  (
    .c({_al_u2514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n205 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n205 ,open_n15123}),
    .q({open_n15127,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [8]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2517|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b8  (
    .c({_al_u2516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n160 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n160 ,open_n15144}),
    .q({open_n15148,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [8]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2518|_al_u2028  (
    .a({open_n15149,_al_u1993_o}),
    .b({_al_u591_o,_al_u591_o}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3:2]),
    .d({_al_u1993_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .f({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }));
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2519|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b8  (
    .c({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n115 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n115 ,open_n15186}),
    .q({open_n15190,\u_cmsdk_mcu/p0_altfunc [8]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2521|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b8  (
    .c({_al_u2520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n70 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n70 ,open_n15207}),
    .q({open_n15211,\u_cmsdk_mcu/p0_outen [8]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u2532|_al_u2533  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/sram_hrdata [10]}),
    .c({\u_cmsdk_mcu/flash_hrdata [10],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]}),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [10],\u_cmsdk_mcu/u_ahb_ram/n13 [10]}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2534|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b2  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,open_n15236}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n275 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n275 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [2]}),
    .q({open_n15252,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2535|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b2  (
    .c({_al_u2476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n238 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n238 ,open_n15269}),
    .q({open_n15273,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [2]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2536|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b2  (
    .c({_al_u2478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n193 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n193 ,open_n15290}),
    .q({open_n15294,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2537|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b2  (
    .c({_al_u2480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n148 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n148 ,open_n15315}),
    .q({open_n15319,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [2]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2538|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b2  (
    .c({_al_u2482_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n103 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n103 ,open_n15340}),
    .q({open_n15344,\u_cmsdk_mcu/p1_altfunc [2]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u2556|_al_u2604  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10]}),
    .c({\u_cmsdk_mcu/flash_hrdata [11],\u_cmsdk_mcu/flash_hrdata [13]}),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [13]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [11],\u_cmsdk_mcu/u_ahb_rom/n13 [13]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2557|_al_u4786  (
    .a({open_n15367,\u_cmsdk_mcu/sram_hrdata [11]}),
    .b({\u_cmsdk_mcu/sram_hrdata [11],\u_cmsdk_mcu/flash_hrdata [11]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [11],_al_u4786_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2558|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b3  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,open_n15390}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n277 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n277 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [3]}),
    .q({open_n15406,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2559|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b3  (
    .c({_al_u2476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n240 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n240 ,open_n15427}),
    .q({open_n15431,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [3]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2560|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b3  (
    .c({_al_u2478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n195 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n195 ,open_n15452}),
    .q({open_n15456,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2561|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b3  (
    .c({_al_u2480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n150 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n150 ,open_n15473}),
    .q({open_n15477,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [3]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2581|_al_u4814  (
    .a({open_n15478,\u_cmsdk_mcu/sram_hrdata [12]}),
    .b({\u_cmsdk_mcu/sram_hrdata [12],\u_cmsdk_mcu/flash_hrdata [12]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [12],_al_u4814_o}));
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2582|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b4  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,open_n15505}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n107 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n279 ,open_n15518}),
    .q({open_n15522,\u_cmsdk_mcu/p0_altfunc [4]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2583|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b4  (
    .c({_al_u2476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n242 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n242 ,open_n15539}),
    .q({open_n15543,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [4]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2584|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b4  (
    .c({_al_u2478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n197 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n197 ,open_n15560}),
    .q({open_n15564,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2605|_al_u4884  (
    .a({open_n15565,\u_cmsdk_mcu/sram_hrdata [13]}),
    .b({\u_cmsdk_mcu/sram_hrdata [13],\u_cmsdk_mcu/flash_hrdata [13]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [13],_al_u4884_o}));
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2606|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b5  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,open_n15588}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n109 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n281 ,open_n15605}),
    .q({open_n15609,\u_cmsdk_mcu/p0_altfunc [5]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2607|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b5  (
    .c({_al_u2476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n244 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n244 ,open_n15626}),
    .q({open_n15630,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [5]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2608|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b5  (
    .c({_al_u2478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n199 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n199 ,open_n15651}),
    .q({open_n15655,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2609|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b5  (
    .c({_al_u2480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n154 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n154 ,open_n15672}),
    .q({open_n15676,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [5]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2629|_al_u4527  (
    .a({open_n15677,\u_cmsdk_mcu/sram_hrdata [14]}),
    .b({\u_cmsdk_mcu/sram_hrdata [14],\u_cmsdk_mcu/flash_hrdata [14]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [14],_al_u4527_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2642|_al_u2985  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 }),
    .b({_al_u2399_o,_al_u2399_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u2642_o,_al_u2985_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(~C*B)))"),
    //.LUT1("(~C*~B*~(~D*~A))"),
    .INIT_LUT0(16'b1010111000000000),
    .INIT_LUT1(16'b0000001100000010),
    .MODE("LOGIC"))
    \_al_u2649|_al_u2648  (
    .a({_al_u2644_o,_al_u682_o}),
    .b({_al_u2646_o,_al_u2647_o}),
    .c({_al_u2648_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u2649_o,_al_u2648_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~B*A)"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(D*C*~B*A)"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2650|_al_u2400  (
    .a({open_n15746,_al_u909_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .d({_al_u2649_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u2650_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B@(A*~(D*~C)))"),
    //.LUTF1("~(B@(A*~(D*~C)))"),
    //.LUTG0("~(B@(A*~(D*~C)))"),
    //.LUTG1("~(B@(A*~(D*~C)))"),
    .INIT_LUTF0(16'b1001001110011001),
    .INIT_LUTF1(16'b1001001110011001),
    .INIT_LUTG0(16'b1001001110011001),
    .INIT_LUTG1(16'b1001001110011001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2651|_al_u2987  (
    .a({_al_u2643_o,_al_u2986_o}),
    .b({_al_u2398_o,_al_u2398_o}),
    .c({_al_u2650_o,_al_u2650_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2664|_al_u4904  (
    .a({open_n15795,\u_cmsdk_mcu/sram_hrdata [15]}),
    .b({\u_cmsdk_mcu/sram_hrdata [15],\u_cmsdk_mcu/flash_hrdata [15]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [15],_al_u4904_o}));
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2665|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b7  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,open_n15818}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n113 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n285 ,open_n15831}),
    .q({open_n15835,\u_cmsdk_mcu/p0_altfunc [7]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u2677|_al_u2706  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]}),
    .c({\u_cmsdk_mcu/flash_hrdata [17],\u_cmsdk_mcu/flash_hrdata [19]}),
    .d({\u_cmsdk_mcu/HWDATA [17],\u_cmsdk_mcu/HWDATA [19]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [17],\u_cmsdk_mcu/u_ahb_rom/n13 [19]}));
  // ../RTL/cmsdk_apb_uart.v(642)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2679|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rxintr_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [1],open_n15860}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable0c ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n117 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n117 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/intr_stat_set [1]}),
    .q({open_n15876,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0]}));  // ../RTL/cmsdk_apb_uart.v(642)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2680|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 ,open_n15879}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n273 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n273 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [1]}),
    .q({open_n15895,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2681|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b1  (
    .c({_al_u2476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n236 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n236 ,open_n15912}),
    .q({open_n15916,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [1]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2682|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b1  (
    .c({_al_u2478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n191 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n191 ,open_n15933}),
    .q({open_n15937,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2683|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b1  (
    .c({_al_u2480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n146 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n146 ,open_n15954}),
    .q({open_n15958,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [1]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2684|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b1  (
    .c({_al_u2482_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n101 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n101 ,open_n15979}),
    .q({open_n15983,\u_cmsdk_mcu/p1_altfunc [1]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2685|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b1  (
    .c({_al_u2484_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n56 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n56 ,open_n16004}),
    .q({open_n16008,\u_cmsdk_mcu/p1_outen [1]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2686|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [1]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n273 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n273 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [1]}),
    .q({open_n16030,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2692|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b9  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n16033}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n289 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n289 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [9]}),
    .q({open_n16053,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2693|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b9  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n252 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n252 ,open_n16074}),
    .q({open_n16078,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [9]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2694|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b9  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n207 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n207 ,open_n16099}),
    .q({open_n16103,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2695|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b9  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n162 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n162 ,open_n16124}),
    .q({open_n16128,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [9]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2696|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b9  (
    .c({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n117 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n117 ,open_n16145}),
    .q({open_n16149,\u_cmsdk_mcu/p1_altfunc [9]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2697|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b9  (
    .c({_al_u2508_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n72 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n72 ,open_n16170}),
    .q({open_n16174,\u_cmsdk_mcu/p1_outen [9]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2698|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b9  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [9]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n289 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n289 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [9]}),
    .q({open_n16196,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2699|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b9  (
    .c({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n252 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n252 ,open_n16217}),
    .q({open_n16221,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [9]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2700|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b9  (
    .c({_al_u2514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n207 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n207 ,open_n16242}),
    .q({open_n16246,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [9]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2701|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b9  (
    .c({_al_u2516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n162 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n162 ,open_n16267}),
    .q({open_n16271,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [9]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2702|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b9  (
    .c({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n117 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n117 ,open_n16288}),
    .q({open_n16292,\u_cmsdk_mcu/p0_altfunc [9]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2703|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b9  (
    .c({_al_u2520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n72 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [9],\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n72 ,open_n16313}),
    .q({open_n16317,\u_cmsdk_mcu/p0_outen [9]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u2704|_al_u3461  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],open_n16320}),
    .c({\u_cmsdk_mcu/flash_hrdata [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({\u_cmsdk_mcu/HWDATA [18],\u_cmsdk_mcu/HWDATA [18]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [18],_al_u3461_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2705|_al_u1835  (
    .a({open_n16341,\u_cmsdk_mcu/sram_hrdata [18]}),
    .b({\u_cmsdk_mcu/sram_hrdata [18],\u_cmsdk_mcu/flash_hrdata [18]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [18],_al_u1835_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2707|_al_u1838  (
    .a({open_n16366,\u_cmsdk_mcu/sram_hrdata [19]}),
    .b({\u_cmsdk_mcu/sram_hrdata [19],\u_cmsdk_mcu/flash_hrdata [19]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [19],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [19],_al_u1838_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2708|_al_u3471  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],open_n16393}),
    .c({\u_cmsdk_mcu/flash_hrdata [20],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({\u_cmsdk_mcu/HWDATA [20],\u_cmsdk_mcu/HWDATA [20]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [20],_al_u3471_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2709|_al_u1841  (
    .a({open_n16418,\u_cmsdk_mcu/sram_hrdata [20]}),
    .b({\u_cmsdk_mcu/sram_hrdata [20],\u_cmsdk_mcu/flash_hrdata [20]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [20],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [20],_al_u1841_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u2710|_al_u2678  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],\u_cmsdk_mcu/sram_hrdata [17]}),
    .c({\u_cmsdk_mcu/flash_hrdata [21],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]}),
    .d({\u_cmsdk_mcu/HWDATA [21],\u_cmsdk_mcu/HWDATA [17]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [21],\u_cmsdk_mcu/u_ahb_ram/n13 [17]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2711|_al_u1843  (
    .a({open_n16465,\u_cmsdk_mcu/sram_hrdata [21]}),
    .b({\u_cmsdk_mcu/sram_hrdata [21],\u_cmsdk_mcu/flash_hrdata [21]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [21],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [21],_al_u1843_o}));
  // ../RTL/cortexm0ds_logic.v(18248)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2716|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6_reg  (
    .a({_al_u2439_o,_al_u1891_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iexow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2272_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n16496,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iexow6 ,_al_u2717_o}),
    .q({open_n16501,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 }));  // ../RTL/cortexm0ds_logic.v(18248)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0011000011111100),
    .MODE("LOGIC"))
    \_al_u2718|_al_u3492  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],open_n16504}),
    .c({\u_cmsdk_mcu/flash_hrdata [24],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({_al_u2717_o,_al_u2717_o}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [24],_al_u3492_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2719|_al_u1850  (
    .a({open_n16525,\u_cmsdk_mcu/sram_hrdata [24]}),
    .b({\u_cmsdk_mcu/sram_hrdata [24],\u_cmsdk_mcu/flash_hrdata [24]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({_al_u2717_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [24],_al_u1850_o}));
  // ../RTL/cortexm0ds_logic.v(18247)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2720|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ,_al_u1971_o}),
    .b({_al_u2261_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awwow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2272_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n16560,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awwow6 ,_al_u2721_o}),
    .q({open_n16565,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 }));  // ../RTL/cortexm0ds_logic.v(18247)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0011000011111100),
    .MODE("LOGIC"))
    \_al_u2722|_al_u3498  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],open_n16568}),
    .c({\u_cmsdk_mcu/flash_hrdata [25],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({_al_u2721_o,_al_u2721_o}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [25],_al_u3498_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"))
    \_al_u2723|_al_u1852  (
    .a({open_n16589,\u_cmsdk_mcu/sram_hrdata [25]}),
    .b({\u_cmsdk_mcu/sram_hrdata [25],\u_cmsdk_mcu/flash_hrdata [25]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({_al_u2721_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [25],_al_u1852_o}));
  // ../RTL/cortexm0ds_logic.v(19947)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(C*~A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2725|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6_reg  (
    .a({_al_u2032_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 }),
    .b({_al_u2455_o,_al_u2272_o}),
    .c({_al_u2724_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n16620,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .f({_al_u2725_o,_al_u2724_o}),
    .q({open_n16625,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 }));  // ../RTL/cortexm0ds_logic.v(19947)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2726|_al_u3503  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],open_n16628}),
    .c({\u_cmsdk_mcu/flash_hrdata [26],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({_al_u2725_o,_al_u2725_o}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [26],_al_u3503_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"))
    \_al_u2727|_al_u1854  (
    .a({open_n16653,\u_cmsdk_mcu/sram_hrdata [26]}),
    .b({\u_cmsdk_mcu/sram_hrdata [26],\u_cmsdk_mcu/flash_hrdata [26]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({_al_u2725_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [26],_al_u1854_o}));
  // ../RTL/cortexm0ds_logic.v(19963)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*~A))"),
    //.LUTF1("(C*~A*~(D*~B))"),
    //.LUTG0("(~(D*C)*~(B*~A))"),
    //.LUTG1("(C*~A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101110111011),
    .INIT_LUTF1(16'b0100000001010000),
    .INIT_LUTG0(16'b0000101110111011),
    .INIT_LUTG1(16'b0100000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2729|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6_reg  (
    .a({_al_u2055_o,_al_u2062_o}),
    .b({_al_u2447_o,_al_u2272_o}),
    .c({_al_u2728_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n16677,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .f({_al_u2729_o,_al_u2728_o}),
    .q({open_n16693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 }));  // ../RTL/cortexm0ds_logic.v(19963)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2731|_al_u1856  (
    .a({open_n16694,\u_cmsdk_mcu/sram_hrdata [27]}),
    .b({\u_cmsdk_mcu/sram_hrdata [27],\u_cmsdk_mcu/flash_hrdata [27]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({_al_u2729_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [27],_al_u1856_o}));
  // ../RTL/cortexm0ds_logic.v(18408)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(B*~A*~(D*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0100000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2733|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6_reg  (
    .a({_al_u2077_o,_al_u2420_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1wow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .c({_al_u2084_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2272_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n16729,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .f({_al_u2733_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1wow6 }),
    .q({open_n16734,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 }));  // ../RTL/cortexm0ds_logic.v(18408)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0011000011111100),
    .MODE("LOGIC"))
    \_al_u2734|_al_u3513  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],open_n16737}),
    .c({\u_cmsdk_mcu/flash_hrdata [28],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({_al_u2733_o,_al_u2733_o}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [28],_al_u3513_o}));
  // ../RTL/cortexm0ds_logic.v(17289)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~A*~(~C*B))"),
    //.LUTF1("(C*~A*~(D*~B))"),
    //.LUTG0("~(~D*~A*~(~C*B))"),
    //.LUTG1("(C*~A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110101110),
    .INIT_LUTF1(16'b0100000001010000),
    .INIT_LUTG0(16'b1111111110101110),
    .INIT_LUTG1(16'b0100000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2741|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6_reg  (
    .a({_al_u2099_o,_al_u2099_o}),
    .b({_al_u2106_o,_al_u1892_o}),
    .c({_al_u2740_o,_al_u2106_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2272_o,_al_u2107_o}),
    .f({_al_u2741_o,\u_cmsdk_mcu/HWDATA [13]}),
    .q({open_n16778,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 }));  // ../RTL/cortexm0ds_logic.v(17289)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .INIT_LUTF0(16'b0011000011111100),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0011000011111100),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2742|_al_u2730  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}),
    .c({\u_cmsdk_mcu/flash_hrdata [29],\u_cmsdk_mcu/flash_hrdata [27]}),
    .d({_al_u2741_o,_al_u2729_o}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [29],\u_cmsdk_mcu/u_ahb_rom/n13 [27]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u2744|_al_u3533  (
    .b({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],open_n16807}),
    .c({\u_cmsdk_mcu/flash_hrdata [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({\u_cmsdk_mcu/HWDATA [16],\u_cmsdk_mcu/HWDATA [16]}),
    .f({\u_cmsdk_mcu/u_ahb_rom/n13 [16],_al_u3533_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2745|_al_u1867  (
    .a({open_n16828,\u_cmsdk_mcu/sram_hrdata [16]}),
    .b({\u_cmsdk_mcu/sram_hrdata [16],\u_cmsdk_mcu/flash_hrdata [16]}),
    .c({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({\u_cmsdk_mcu/HWDATA [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n13 [16],_al_u1867_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~A*~(~B*~(D*~C)))"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~A*~(~B*~(D*~C)))"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0100010101000100),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0100010101000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2746|_al_u916  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 }),
    .f({_al_u2746_o,_al_u916_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~B*~(~D*C*A))"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0011001100010011),
    .MODE("LOGIC"))
    \_al_u2747|_al_u1383  (
    .a({_al_u916_o,open_n16877}),
    .b({_al_u2746_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,_al_u916_o}),
    .f({_al_u2747_o,_al_u1383_o}));
  // ../RTL/cortexm0ds_logic.v(17657)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~B*D)"),
    //.LUT1("(B*~(C*~(D*A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111111111),
    .INIT_LUT1(16'b1000110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2748|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6_reg  (
    .a({_al_u1765_o,open_n16898}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ,_al_u2748_o}),
    .c({_al_u2747_o,_al_u2751_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 }),
    .f({_al_u2748_o,open_n16912}),
    .q({open_n16916,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 }));  // ../RTL/cortexm0ds_logic.v(17657)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u2750|_al_u912  (
    .b({_al_u2749_o,open_n16919}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({_al_u912_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv }),
    .f({_al_u2750_o,_al_u912_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2751|_al_u918  (
    .a({open_n16940,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv ,_al_u916_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K75iu6_lutinv }),
    .d({_al_u2750_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .f({_al_u2751_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aj1ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("(~C*~A*~(~D*B))"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("(~C*~A*~(~D*B))"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000010100000001),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b0000010100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2756|_al_u2755  (
    .a({_al_u2754_o,_al_u2365_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({_al_u2755_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u2756_o,_al_u2755_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2758|_al_u1805  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u2758_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*A*~(D*~B))"),
    //.LUTF1("(~D*~A*~(C*B))"),
    //.LUTG0("(~C*A*~(D*~B))"),
    //.LUTG1("(~D*~A*~(C*B))"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000000000010101),
    .INIT_LUTG0(16'b0000100000001010),
    .INIT_LUTG1(16'b0000000000010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2760|_al_u2759  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ,_al_u903_o}),
    .b({_al_u681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .c({_al_u2758_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u2759_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u2760_o,_al_u2759_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(~C*B)))"),
    //.LUT1("(C*A*~(D*B))"),
    .INIT_LUT0(16'b1010111000000000),
    .INIT_LUT1(16'b0010000010100000),
    .MODE("LOGIC"))
    \_al_u2761|_al_u2757  (
    .a({_al_u2756_o,_al_u1782_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .c({_al_u2760_o,_al_u1271_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .f({_al_u2761_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2763|_al_u2762  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({_al_u2365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u2763_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2765|_al_u2764  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({_al_u2764_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ,_al_u2764_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"))
    \_al_u2766|_al_u2832  (
    .a({_al_u2763_o,open_n17113}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv }),
    .f({_al_u2766_o,_al_u2832_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B*A))"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~D*~(~C*~B*A))"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0000000011111101),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000000011111101),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2768|_al_u3687  (
    .a({open_n17134,_al_u2767_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ,_al_u2369_o}),
    .c({_al_u2767_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Io9ow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~A*~(~D*B)))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*~(~A*~(~D*B)))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1010000011100000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1010000011100000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2769|_al_u3858  (
    .a({open_n17159,_al_u2766_o}),
    .b({open_n17160,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({_al_u2766_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ,_al_u3858_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2771|_al_u2770  (
    .c({_al_u2770_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .f({_al_u2771_o,_al_u2770_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(A*~(~B*~(D*~C)))"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b1000101010001000),
    .MODE("LOGIC"))
    \_al_u2773|_al_u2772  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,open_n17209}),
    .b({_al_u2772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({_al_u2770_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv }),
    .f({_al_u2773_o,_al_u2772_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~B*~(D*C*A))"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0001001100110011),
    .MODE("LOGIC"))
    \_al_u2776|_al_u2774  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,open_n17230}),
    .b({_al_u2774_o,_al_u909_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u2776_o,_al_u2774_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~(~D*A))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*~B*~(~D*A))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .INIT_LUTF0(16'b0011000000010000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2778|_al_u2777  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv ,_al_u2771_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ,_al_u2773_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,_al_u2776_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u2778_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2779|_al_u1346  (
    .b({_al_u1346_o,open_n17277}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u2779_o,_al_u1346_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u277|_al_u283  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u2780|_al_u1264  (
    .b({_al_u1264_o,open_n17332}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u2779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 ,_al_u1264_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2782|_al_u2781  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u2782_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0000001010100010),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0000001010100010),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2783|_al_u3407  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3kiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u2782_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u2783_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 }));
  // ../RTL/cortexm0ds_logic.v(18707)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(B*A*~(~D*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b1000100010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2784|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6_reg  (
    .a({_al_u2761_o,open_n17405}),
    .b({_al_u2778_o,open_n17406}),
    .c({_al_u2783_o,_al_u2791_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ,_al_u2784_o}),
    .f({_al_u2784_o,open_n17420}),
    .q({open_n17424,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 }));  // ../RTL/cortexm0ds_logic.v(18707)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D@C@B@A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0110100110010110),
    .MODE("LOGIC"))
    \_al_u2785|_al_u2380  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .f({_al_u2785_o,_al_u2380_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*C))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2787|_al_u4339  (
    .a({open_n17445,_al_u4325_o}),
    .b({open_n17446,_al_u4338_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,_al_u3608_o}),
    .d({_al_u2786_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({_al_u2787_o,_al_u4339_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2788|_al_u3311  (
    .b({open_n17469,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({_al_u2787_o,_al_u2787_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2789|_al_u1356  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,open_n17494}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ,open_n17495}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u2789_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u278|_al_u282  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B*~A))"),
    //.LUT1("(C*B*~D)"),
    .INIT_LUT0(16'b0000000011111110),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"))
    \_al_u2794|_al_u2795  (
    .a({open_n17548,_al_u2794_o}),
    .b({_al_u2793_o,_al_u1643_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ,_al_u1777_o}),
    .d({_al_u1906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({_al_u2794_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkliu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2796|_al_u7208  (
    .b({open_n17571,_al_u1299_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 }),
    .d({_al_u1906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ,_al_u7208_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2798|_al_u609  (
    .c({_al_u609_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u1788_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ,_al_u609_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u279|_al_u281  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [5]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B@D))"),
    //.LUTF1("(~D*~C*~(B*A))"),
    //.LUTG0("(~C*(B@D))"),
    //.LUTG1("(~D*~C*~(B*A))"),
    .INIT_LUTF0(16'b0000001100001100),
    .INIT_LUTF1(16'b0000000000000111),
    .INIT_LUTG0(16'b0000001100001100),
    .INIT_LUTG1(16'b0000000000000111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2803|_al_u2802  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ,open_n17648}),
    .b({_al_u1658_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({_al_u1817_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u2802_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u2803_o,_al_u2802_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*B*~A))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(C*~(D*B*~A))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b1011000011110000),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011000011110000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2804|_al_u2800  (
    .a({_al_u2800_o,_al_u1336_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .c({_al_u2803_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u2804_o,_al_u2800_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*~A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*~A))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0010101000111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0010101000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2805|_al_u932  (
    .a({_al_u2804_o,open_n17697}),
    .b({_al_u932_o,open_n17698}),
    .c({_al_u2403_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ,_al_u932_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2808|_al_u2807  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ,open_n17725}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u1342_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u2808_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B))"),
    //.LUTF1("(~B*A*~(~D*~C))"),
    //.LUTG0("(D*~(C*~B))"),
    //.LUTG1("(~B*A*~(~D*~C))"),
    .INIT_LUTF0(16'b1100111100000000),
    .INIT_LUTF1(16'b0010001000100000),
    .INIT_LUTG0(16'b1100111100000000),
    .INIT_LUTG1(16'b0010001000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2810|_al_u2809  (
    .a({_al_u2808_o,open_n17750}),
    .b({_al_u2809_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u1658_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .f({_al_u2810_o,_al_u2809_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2814|_al_u2813  (
    .a({_al_u2810_o,open_n17775}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 ,open_n17776}),
    .c({_al_u932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u2813_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ,_al_u2813_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~(B*~A))"),
    //.LUTF1("(C*~(~B*~D))"),
    //.LUTG0("(~D*C*~(B*~A))"),
    //.LUTG1("(C*~(~B*~D))"),
    .INIT_LUTF0(16'b0000000010110000),
    .INIT_LUTF1(16'b1111000011000000),
    .INIT_LUTG0(16'b0000000010110000),
    .INIT_LUTG1(16'b1111000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2816|_al_u2815  (
    .a({open_n17801,_al_u607_o}),
    .b({_al_u2387_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u2815_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u2816_o,_al_u2815_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(~A*~(~D*B)))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(~A*~(~D*B)))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010000011100000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010000011100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2817|_al_u682  (
    .a({_al_u682_o,open_n17826}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ,open_n17827}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u2817_o,_al_u682_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*D))"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(~C*~(B*D))"),
    //.LUTG1("(~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000001100001111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001100001111),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2819|_al_u2820  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ,open_n17852}),
    .b({_al_u2816_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 }),
    .c({_al_u2817_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u2818_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2822|_al_u2821  (
    .b({open_n17879,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({_al_u2365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b0100010001010000),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u2824|_al_u2823  (
    .a({open_n17900,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .b({_al_u2772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u2824_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000001100001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2826|_al_u1370  (
    .b({open_n17923,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ,_al_u1370_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(A*~(B*~(D*~C)))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(A*~(B*~(D*~C)))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0010101000100010),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0010101000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2827|_al_u2835  (
    .a({_al_u2825_o,open_n17944}),
    .b({_al_u2771_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,_al_u2771_o}),
    .f({_al_u2827_o,_al_u2835_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*~C))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1000000010001000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2828|_al_u3843  (
    .a({open_n17969,_al_u2361_o}),
    .b({open_n17970,_al_u3840_o}),
    .c({_al_u2772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,_al_u2764_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 ,_al_u3843_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2830|_al_u2829  (
    .b({_al_u2829_o,open_n17993}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 ,_al_u2829_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u2831|_al_u6253  (
    .a({open_n18014,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 ,_al_u1812_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mldpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ,_al_u6253_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u2833|_al_u3421  (
    .a({open_n18035,_al_u3420_o}),
    .b({_al_u2832_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmiiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8iiu6 ,_al_u3421_o}));
  // ../RTL/cortexm0ds_logic.v(18701)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2834|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K8iiu6 ,_al_u2841_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2827_o,_al_u2834_o}),
    .f({_al_u2834_o,open_n18071}),
    .q({open_n18075,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 }));  // ../RTL/cortexm0ds_logic.v(18701)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(D*~C)))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0100110001000100),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u2838|_al_u2837  (
    .a({open_n18076,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .b({_al_u2836_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .c({_al_u2837_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u2771_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ,_al_u2837_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2840|_al_u2839  (
    .b({_al_u2373_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .c({_al_u2770_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({_al_u2839_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u2840_o,_al_u2839_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~D*~C*B*~A)"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("LOGIC"))
    \_al_u2841|_al_u3608  (
    .a({_al_u2835_o,_al_u2835_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 }),
    .c({_al_u2763_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u2840_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u2841_o,_al_u3608_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u2843|_al_u2811  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ,open_n18145}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u2843_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*~A)"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~D*~C*B*~A)"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2845|_al_u3661  (
    .a({open_n18166,_al_u1643_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u2845_o,_al_u3661_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2847|_al_u3104  (
    .a({open_n18191,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .b({open_n18192,_al_u932_o}),
    .c({_al_u1346_o,_al_u1346_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }),
    .f({_al_u2847_o,_al_u3104_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2848|_al_u5982  (
    .b({open_n18219,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 }),
    .c({_al_u2847_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .d({_al_u2846_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk5ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u2849|_al_u1332  (
    .a({open_n18244,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u2849_o,_al_u1332_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~(B*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~D*~C*~(B*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000000000111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000000111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2850|_al_u2858  (
    .a({open_n18265,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 }),
    .b({_al_u1336_o,_al_u1812_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u2849_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ,_al_u2858_o}));
  // ../RTL/cortexm0ds_logic.v(17500)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2851|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6_reg  (
    .a({open_n18290,_al_u4488_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ja5iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv ,open_n18304}),
    .q({open_n18308,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 }));  // ../RTL/cortexm0ds_logic.v(17500)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2853|_al_u3891  (
    .b({open_n18311,_al_u3624_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ,_al_u3891_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2854|_al_u2818  (
    .b({open_n18338,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u1583_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ,_al_u2818_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(~A*~(~D*~(~C*~B)))"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b0101010100000001),
    .MODE("LOGIC"))
    \_al_u2855|_al_u3570  (
    .a({_al_u2847_o,open_n18359}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv }),
    .f({_al_u2855_o,_al_u3570_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~(~B*~D))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000011000000),
    .MODE("LOGIC"))
    \_al_u2856|_al_u675  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ,open_n18382}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn ,\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn }),
    .d({_al_u1385_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17506)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(D*~(C*~B*A))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1101111100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2857|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbopw6_reg  (
    .a({open_n18403,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv }),
    .b({open_n18404,_al_u2857_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ,_al_u2858_o}),
    .clk(XTAL1_wire),
    .d({_al_u2855_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2857_o,open_n18422}),
    .q({open_n18426,\u_cmsdk_mcu/u_cmsdk_mcu_system/SLEEPHOLDACKn }));  // ../RTL/cortexm0ds_logic.v(17506)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u2861|_al_u1344  (
    .a({_al_u1344_o,open_n18427}),
    .b({_al_u2403_o,open_n18428}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u2861_o,_al_u1344_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(B*~(D*C*A))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(B*~(D*C*A))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0100110011001100),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2863|_al_u1340  (
    .a({_al_u2860_o,open_n18449}),
    .b({_al_u2862_o,open_n18450}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u2863_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2864|_al_u2865  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .c({_al_u2770_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 ,_al_u2865_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~D*B*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2866|_al_u3123  (
    .a({open_n18499,_al_u2866_o}),
    .b({open_n18500,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,_al_u3122_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u2866_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~(~D*B)*~(C*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0101111100010011),
    .MODE("LOGIC"))
    \_al_u2867|_al_u679  (
    .a({_al_u1806_o,open_n18521}),
    .b({_al_u2866_o,open_n18522}),
    .c({_al_u679_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u2867_o,_al_u679_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(~A*~(D*C)))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1100100010001000),
    .MODE("LOGIC"))
    \_al_u2869|_al_u2868  (
    .a({_al_u1812_o,open_n18543}),
    .b({_al_u2868_o,open_n18544}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .f({_al_u2869_o,_al_u2868_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~(~D*B)*~(C*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0101111100010011),
    .MODE("LOGIC"))
    \_al_u2870|_al_u1907  (
    .a({_al_u609_o,open_n18565}),
    .b({_al_u1346_o,open_n18566}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u1907_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u2870_o,_al_u1907_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(D*~C)))"),
    //.LUT1("(D*~C*~(~B*A))"),
    .INIT_LUT0(16'b0010101000100010),
    .INIT_LUT1(16'b0000110100000000),
    .MODE("LOGIC"))
    \_al_u2872|_al_u2871  (
    .a({_al_u1643_o,_al_u2870_o}),
    .b({_al_u2867_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({_al_u2869_o,_al_u1266_o}),
    .d({_al_u2871_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u2872_o,_al_u2871_o}));
  // ../RTL/cortexm0ds_logic.v(17759)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C*~B*~(~D*~A))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C*~B*~(~D*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110100010001),
    .INIT_LUTF1(16'b0011000000100000),
    .INIT_LUTG0(16'b1111110100010001),
    .INIT_LUTG1(16'b0011000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2873|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6_reg  (
    .a({_al_u2863_o,_al_u2873_o}),
    .b({_al_u2865_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({_al_u2872_o,_al_u1817_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2873_o,open_n18624}),
    .q({open_n18628,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }));  // ../RTL/cortexm0ds_logic.v(17759)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(B@(D*~(C*~A)))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(B@(D*~(C*~A)))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1001110000110011),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1001110000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2876|_al_u2875  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ,_al_u2399_o}),
    .b({_al_u2398_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 }),
    .c({_al_u2412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 }),
    .d({_al_u2875_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10],_al_u2875_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u2878|_al_u2877  (
    .a({open_n18653,_al_u2399_o}),
    .b({_al_u2877_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kc6ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({_al_u2878_o,_al_u2877_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2881|_al_u2880  (
    .a({open_n18674,_al_u2849_o}),
    .b({open_n18675,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .d({_al_u2650_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u2881_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef7ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B@(A*~(D*~C)))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("~(B@(A*~(D*~C)))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .INIT_LUTF0(16'b1001001110011001),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1001001110011001),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2882|_al_u3036  (
    .a({_al_u1882_o,_al_u3035_o}),
    .b({_al_u2881_o,_al_u2398_o}),
    .c({_al_u2412_o,_al_u2881_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }),
    .f({_al_u2882_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B))"),
    //.LUTF1("~(C@D)"),
    //.LUTG0("(D*~(C*~B))"),
    //.LUTG1("~(C@D)"),
    .INIT_LUTF0(16'b1100111100000000),
    .INIT_LUTF1(16'b1111000000001111),
    .INIT_LUTG0(16'b1100111100000000),
    .INIT_LUTG1(16'b1111000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2883|_al_u2643  (
    .b({open_n18722,_al_u1952_o}),
    .c({_al_u2398_o,_al_u2412_o}),
    .d({_al_u2882_o,_al_u2642_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0],_al_u2643_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2884|_al_u2890  (
    .c({_al_u588_o,_al_u591_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2886|_al_u2888  (
    .c({_al_u593_o,_al_u585_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 }));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2892|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b10  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n18801}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [10]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n291 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n291 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [10]}),
    .q({open_n18821,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2893|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b10  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n254 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n254 ,open_n18838}),
    .q({open_n18842,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [10]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2894|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b10  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n209 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n209 ,open_n18859}),
    .q({open_n18863,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2895|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b10  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n164 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n164 ,open_n18884}),
    .q({open_n18888,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [10]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2896|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b10  (
    .c({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n119 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n119 ,open_n18905}),
    .q({open_n18909,\u_cmsdk_mcu/p1_altfunc [10]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2897|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b10  (
    .c({_al_u2508_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n74 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n74 ,open_n18930}),
    .q({open_n18934,\u_cmsdk_mcu/p1_outen [10]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2898|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b10  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [10]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [10]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n291 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n291 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [10]}),
    .q({open_n18952,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2899|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b10  (
    .c({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n254 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n254 ,open_n18969}),
    .q({open_n18973,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [10]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2900|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b10  (
    .c({_al_u2514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n209 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n209 ,open_n18990}),
    .q({open_n18994,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [10]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2901|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b10  (
    .c({_al_u2516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n164 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n164 ,open_n19015}),
    .q({open_n19019,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [10]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2902|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b10  (
    .c({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n119 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n119 ,open_n19040}),
    .q({open_n19044,\u_cmsdk_mcu/p0_altfunc [10]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2903|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b10  (
    .c({_al_u2520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n74 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [10],\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n74 ,open_n19065}),
    .q({open_n19069,\u_cmsdk_mcu/p0_outen [10]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2906|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b11  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n19072}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [11]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n293 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n293 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [11]}),
    .q({open_n19092,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2907|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b11  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n256 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n256 ,open_n19109}),
    .q({open_n19113,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [11]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2908|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b11  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n211 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n211 ,open_n19130}),
    .q({open_n19134,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2909|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b11  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n166 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n166 ,open_n19151}),
    .q({open_n19155,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [11]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2910|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b11  (
    .c({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n121 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n121 ,open_n19176}),
    .q({open_n19180,\u_cmsdk_mcu/p1_altfunc [11]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2911|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b11  (
    .c({_al_u2508_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n76 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n76 ,open_n19197}),
    .q({open_n19201,\u_cmsdk_mcu/p1_outen [11]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2912|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b11  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [11]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [11]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n293 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n293 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [11]}),
    .q({open_n19223,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2913|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b11  (
    .c({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n256 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n256 ,open_n19240}),
    .q({open_n19244,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [11]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2914|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b11  (
    .c({_al_u2514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n211 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n211 ,open_n19261}),
    .q({open_n19265,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [11]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2915|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b11  (
    .c({_al_u2516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n166 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n166 ,open_n19282}),
    .q({open_n19286,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [11]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2916|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b11  (
    .c({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n121 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n121 ,open_n19307}),
    .q({open_n19311,\u_cmsdk_mcu/p0_altfunc [11]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2917|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b11  (
    .c({_al_u2520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n76 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n76 ,open_n19328}),
    .q({open_n19332,\u_cmsdk_mcu/p0_outen [11]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("~(B@(D*~(C*~A)))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1001110000110011),
    .MODE("LOGIC"))
    \_al_u2922|_al_u2921  (
    .a({_al_u2062_o,open_n19333}),
    .b({_al_u2398_o,_al_u2399_o}),
    .c({_al_u2412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({_al_u2921_o,_al_u2920_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 ,_al_u2921_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2923|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b12  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n19356}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [12]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n295 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n295 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [12]}),
    .q({open_n19372,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2924|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b12  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n258 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n258 ,open_n19393}),
    .q({open_n19397,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [12]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2925|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b12  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n213 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n213 ,open_n19414}),
    .q({open_n19418,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2926|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b12  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n168 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n168 ,open_n19439}),
    .q({open_n19443,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [12]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2927|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b12  (
    .c({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n123 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n123 ,open_n19464}),
    .q({open_n19468,\u_cmsdk_mcu/p1_altfunc [12]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2928|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b12  (
    .c({_al_u2508_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n78 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n78 ,open_n19485}),
    .q({open_n19489,\u_cmsdk_mcu/p1_outen [12]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2929|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b12  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [12]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [12]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n295 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n295 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [12]}),
    .q({open_n19511,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2930|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b12  (
    .c({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n258 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n258 ,open_n19528}),
    .q({open_n19532,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [12]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2931|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b12  (
    .c({_al_u2514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n213 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n213 ,open_n19553}),
    .q({open_n19557,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [12]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2932|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b12  (
    .c({_al_u2516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n168 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n168 ,open_n19578}),
    .q({open_n19582,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [12]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2933|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b12  (
    .c({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n123 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n123 ,open_n19603}),
    .q({open_n19607,\u_cmsdk_mcu/p0_altfunc [12]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2934|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b12  (
    .c({_al_u2520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n78 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n78 ,open_n19624}),
    .q({open_n19628,\u_cmsdk_mcu/p0_outen [12]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("~(B@(D*~(C*~A)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1001110000110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u2937|_al_u2938  (
    .a({open_n19629,_al_u2084_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u2937_o}),
    .f({_al_u2937_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 }));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2939|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b13  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n19652}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [13]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n297 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n297 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [13]}),
    .q({open_n19668,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2940|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b13  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n260 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n260 ,open_n19685}),
    .q({open_n19689,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [13]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2941|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b13  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n215 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n215 ,open_n19706}),
    .q({open_n19710,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2942|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b13  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n170 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n170 ,open_n19727}),
    .q({open_n19731,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [13]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2943|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b13  (
    .c({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n125 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n125 ,open_n19752}),
    .q({open_n19756,\u_cmsdk_mcu/p1_altfunc [13]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2944|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b13  (
    .c({_al_u2508_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n80 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n80 ,open_n19773}),
    .q({open_n19777,\u_cmsdk_mcu/p1_outen [13]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2945|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b13  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [13]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [13]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n297 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n297 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [13]}),
    .q({open_n19795,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2946|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b13  (
    .c({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n260 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n260 ,open_n19812}),
    .q({open_n19816,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [13]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2947|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b13  (
    .c({_al_u2514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n215 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n215 ,open_n19833}),
    .q({open_n19837,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [13]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2948|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b13  (
    .c({_al_u2516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n170 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n170 ,open_n19854}),
    .q({open_n19858,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [13]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2949|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b13  (
    .c({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n125 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n125 ,open_n19879}),
    .q({open_n19883,\u_cmsdk_mcu/p0_altfunc [13]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u294|_al_u4657  (
    .c({\u_cmsdk_mcu/u_ahb_ram/we ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0]}),
    .d({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [12],_al_u4603_o}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n16 ,_al_u4657_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2950|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b13  (
    .c({_al_u2520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n80 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n80 ,open_n19928}),
    .q({open_n19932,\u_cmsdk_mcu/p0_outen [13]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B@(D*~(C*~A)))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B@(D*~(C*~A)))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1001110000110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1001110000110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2953|_al_u2954  (
    .a({open_n19933,_al_u2106_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u2953_o}),
    .f({_al_u2953_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 }));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2955|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b14  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n19960}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [14]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n299 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n299 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [14]}),
    .q({open_n19980,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2956|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b14  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n262 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [14],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n262 ,open_n20001}),
    .q({open_n20005,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [14]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2957|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b14  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n217 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [14],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n217 ,open_n20022}),
    .q({open_n20026,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2958|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b14  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n172 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [14],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n172 ,open_n20043}),
    .q({open_n20047,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [14]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B@(D*~(C*~A)))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B@(D*~(C*~A)))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1001110000110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1001110000110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2969|_al_u2970  (
    .a({open_n20048,_al_u2128_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u2969_o}),
    .f({_al_u2969_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 }));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2971|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b15  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write1 ,open_n20075}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [15]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n301 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n301 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [15]}),
    .q({open_n20095,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2972|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b15  (
    .c({_al_u2500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n264 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n264 ,open_n20116}),
    .q({open_n20120,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [15]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2973|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b15  (
    .c({_al_u2502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n219 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n219 ,open_n20141}),
    .q({open_n20145,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2974|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b15  (
    .c({_al_u2504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n174 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n174 ,open_n20166}),
    .q({open_n20170,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [15]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2975|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b15  (
    .c({_al_u2506_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n129 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n129 ,open_n20187}),
    .q({open_n20191,\u_cmsdk_mcu/p1_altfunc [15]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2976|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b15  (
    .c({_al_u2508_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n84 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n84 ,open_n20212}),
    .q({open_n20216,\u_cmsdk_mcu/p1_outen [15]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("~(~C*~(B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111110011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2977|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b15  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [15]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [15]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n301 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n301 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [15]}),
    .q({open_n20238,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2978|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b15  (
    .c({_al_u2512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n264 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n264 ,open_n20259}),
    .q({open_n20263,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [15]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2979|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b15  (
    .c({_al_u2514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n219 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n219 ,open_n20284}),
    .q({open_n20288,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [15]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2980|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg4_b15  (
    .c({_al_u2516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n136 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n174 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n174 ,open_n20309}),
    .q({open_n20313,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [15]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2981|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg3_b15  (
    .c({_al_u2518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n91 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n129 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n129 ,open_n20330}),
    .q({open_n20334,\u_cmsdk_mcu/p0_altfunc [15]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2982|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b15  (
    .c({_al_u2520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n84 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [15],\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n84 ,open_n20355}),
    .q({open_n20359,\u_cmsdk_mcu/p0_outen [15]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cortexm0ds_logic.v(19665)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(D*~(C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2986|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6_reg  (
    .b({_al_u1961_o,_al_u1961_o}),
    .c({_al_u2412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2985_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxow6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2986_o,\u_cmsdk_mcu/HWDATA [23]}),
    .q({open_n20377,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 }));  // ../RTL/cortexm0ds_logic.v(19665)
  EG_PHY_MSLICE #(
    //.LUT0("~(B@(D*~(C*~A)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1001110000110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u2988|_al_u2989  (
    .a({open_n20378,_al_u2150_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u2988_o}),
    .f({_al_u2988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(B@(D*~(C*~A)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1001110000110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u2990|_al_u2991  (
    .a({open_n20399,_al_u2171_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u2990_o}),
    .f({_al_u2990_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 }));
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(~C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2992|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b4  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .clk(XTAL1_wire),
    .d({_al_u497_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}),
    .mi({open_n20432,\u_cmsdk_mcu/HADDR [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u2992_o,_al_u498_o}),
    .q({open_n20436,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6]}));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2994|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe [0],open_n20439}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable ,\u_cmsdk_mcu/HWRITE }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ,open_n20452}),
    .q({open_n20456,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable }));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  // ../RTL/cmsdk_apb_uart.v(368)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111111111111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u299|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated_reg  (
    .b({uart0_txen_pad,open_n20459}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n46 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 }),
    .q({open_n20475,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated }));  // ../RTL/cmsdk_apb_uart.v(368)
  EG_PHY_MSLICE #(
    //.LUT0("~(B@(D*~(C*~A)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1001110000110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3000|_al_u3001  (
    .a({open_n20476,_al_u2208_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u3000_o}),
    .f({_al_u3000_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B@(D*~(C*~A)))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B@(D*~(C*~A)))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1001110000110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1001110000110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3002|_al_u3003  (
    .a({open_n20497,_al_u2217_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u3002_o}),
    .f({_al_u3002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B@(D*~(C*~A)))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B@(D*~(C*~A)))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1001110000110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1001110000110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3004|_al_u3005  (
    .a({open_n20522,_al_u2225_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u3004_o}),
    .f({_al_u3004_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(B@(D*~(C*~A)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1001110000110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3006|_al_u3007  (
    .a({open_n20547,_al_u2235_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u3006_o}),
    .f({_al_u3006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 }));
  // ../RTL/cortexm0ds_logic.v(20093)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(B@(D*~(C*~A)))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(B@(D*~(C*~A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b1001110000110011),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b1001110000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3009|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6_reg  (
    .a({_al_u2244_o,open_n20568}),
    .b({_al_u2398_o,_al_u2244_o}),
    .c({_al_u2412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u3008_o,_al_u2237_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ,\u_cmsdk_mcu/HWDATA [22]}),
    .q({open_n20588,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 }));  // ../RTL/cortexm0ds_logic.v(20093)
  // ../RTL/cortexm0ds_logic.v(18417)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u300|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ,open_n20605}),
    .q({open_n20609,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 }));  // ../RTL/cortexm0ds_logic.v(18417)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUTF1("~(B@(D*~(C*~A)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUTG1("~(B@(D*~(C*~A)))"),
    .INIT_LUTF0(16'b0001001111110101),
    .INIT_LUTF1(16'b1001110000110011),
    .INIT_LUTG0(16'b0001001111110101),
    .INIT_LUTG1(16'b1001110000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3011|_al_u3010  (
    .a({_al_u2252_o,_al_u2399_o}),
    .b({_al_u2398_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 }),
    .c({_al_u2412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({_al_u3010_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23],_al_u3010_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B@(D*~(C*~A)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1001110000110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3012|_al_u3013  (
    .a({open_n20634,_al_u2289_o}),
    .b({_al_u2399_o,_al_u2398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ,_al_u2412_o}),
    .d({_al_u2920_o,_al_u3012_o}),
    .f({_al_u3012_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3015|_al_u3014  (
    .b({open_n20657,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv ,_al_u607_o}),
    .f({_al_u3015_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(D*C)*~(B*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(D*C)*~(B*A))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000011101110111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3020|_al_u3019  (
    .a({_al_u1342_o,open_n20682}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ,open_n20683}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u3020_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUT1("(B*~(D*~C*~A))"),
    .INIT_LUT0(16'b0000110011111100),
    .INIT_LUT1(16'b1100100011001100),
    .MODE("LOGIC"))
    \_al_u3021|_al_u3017  (
    .a({_al_u3017_o,open_n20708}),
    .b({_al_u3020_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 }),
    .f({_al_u3021_o,_al_u3017_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"))
    \_al_u3023|_al_u5993  (
    .a({_al_u1943_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwzhu6 }),
    .b({_al_u3022_o,_al_u607_o}),
    .c({_al_u2412_o,_al_u932_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 }),
    .f({_al_u3023_o,_al_u5993_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("~(B@(C*D))"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1100001100110011),
    .MODE("LOGIC"))
    \_al_u3025|_al_u3024  (
    .a({open_n20749,_al_u2650_o}),
    .b({_al_u2398_o,_al_u2399_o}),
    .c({_al_u3024_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 }),
    .d({_al_u3023_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5],_al_u3024_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3026|_al_u3029  (
    .a({_al_u1925_o,_al_u1934_o}),
    .b({_al_u3022_o,_al_u3022_o}),
    .c({_al_u2412_o,_al_u2412_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }),
    .f({_al_u3026_o,_al_u3029_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*~A))"),
    //.LUTF1("~(B@(C*D))"),
    //.LUTG0("(~(C*B)*~(D*~A))"),
    //.LUTG1("~(B@(C*D))"),
    .INIT_LUTF0(16'b0010101000111111),
    .INIT_LUTF1(16'b1100001100110011),
    .INIT_LUTG0(16'b0010101000111111),
    .INIT_LUTG1(16'b1100001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3028|_al_u3027  (
    .a({open_n20794,_al_u2650_o}),
    .b({_al_u2398_o,_al_u2399_o}),
    .c({_al_u3027_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .d({_al_u3026_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3],_al_u3027_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("~(B@(C*D))"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1100001100110011),
    .MODE("LOGIC"))
    \_al_u3031|_al_u3030  (
    .a({open_n20819,_al_u2650_o}),
    .b({_al_u2398_o,_al_u2399_o}),
    .c({_al_u3030_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .d({_al_u3029_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [4],_al_u3030_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("~(B@(A*~(D*~C)))"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b1001001110011001),
    .MODE("LOGIC"))
    \_al_u3033|_al_u3032  (
    .a({_al_u3032_o,_al_u1968_o}),
    .b({_al_u2398_o,_al_u2412_o}),
    .c({_al_u2881_o,_al_u2399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1],_al_u3032_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u3035|_al_u3034  (
    .a({open_n20860,_al_u3022_o}),
    .b({_al_u1916_o,_al_u2399_o}),
    .c({_al_u2412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .d({_al_u3034_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 }),
    .f({_al_u3035_o,_al_u3034_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3039|_al_u3038  (
    .a({open_n20881,_al_u1048_o}),
    .b({open_n20882,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n12_lutinv }));
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~(D*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000100000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3041|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b2  (
    .a({\u_cmsdk_mcu/HWDATA [0],open_n20903}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 ,open_n20904}),
    .c({_al_u3040_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [0],_al_u3047_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3041_o,open_n20918}),
    .q({open_n20922,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [2]}));  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~C*~B*~(D*A))"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000000100000011),
    .MODE("LOGIC"))
    \_al_u3079|_al_u3078  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ,_al_u695_o}),
    .b({_al_u3078_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({_al_u1264_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u2371_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3079_o,_al_u3078_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3081|_al_u3207  (
    .c({_al_u2376_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv }),
    .f({_al_u3081_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*~(D*B*~A))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000101100001111),
    .MODE("LOGIC"))
    \_al_u3083|_al_u3082  (
    .a({_al_u1812_o,open_n20971}),
    .b({_al_u1799_o,_al_u2813_o}),
    .c({_al_u3082_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,_al_u604_o}),
    .f({_al_u3083_o,_al_u3082_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~(~B*~A))"),
    //.LUT1("(C*~B*~(~D*A))"),
    .INIT_LUT0(16'b1110000000000000),
    .INIT_LUT1(16'b0011000000010000),
    .MODE("LOGIC"))
    \_al_u3084|_al_u4036  (
    .a({_al_u1801_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 }),
    .b({_al_u3081_o,_al_u3081_o}),
    .c({_al_u3083_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ,_al_u4036_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3085|_al_u1801  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 }),
    .f({_al_u3085_o,_al_u1801_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*B)*~(~D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b1111001101010001),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u3087|_al_u3086  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 }),
    .b({_al_u3086_o,_al_u3085_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3087_o,_al_u3086_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3089|_al_u3088  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ,open_n21062}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u1802_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*~C*B))"),
    //.LUT1("(B*~(A*~(D*C)))"),
    .INIT_LUT0(16'b0101000101010101),
    .INIT_LUT1(16'b1100010001000100),
    .MODE("LOGIC"))
    \_al_u3092|_al_u3091  (
    .a({_al_u3091_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjiow6 }),
    .b({_al_u2361_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({_al_u2365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3092_o,_al_u3091_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~C*B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~(~D*~C*B))"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b1010101010100010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1010101010100010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3093|_al_u3080  (
    .a({_al_u3080_o,_al_u3079_o}),
    .b({_al_u3087_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u3092_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 ,_al_u3080_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3094|_al_u7153  (
    .a({open_n21131,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 ,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [2]}),
    .f({_al_u3094_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwgow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3099|_al_u3100  (
    .a({open_n21156,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkjiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njjiu6_lutinv }),
    .d({_al_u1812_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Njjiu6_lutinv ,_al_u3100_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3101|_al_u1665  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ,open_n21183}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u3101_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3102|_al_u1324  (
    .b({_al_u2758_o,open_n21206}),
    .c({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u3101_o,_al_u1266_o}),
    .f({_al_u3102_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3105|_al_u3103  (
    .b({_al_u3104_o,open_n21229}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u3103_o,_al_u1266_o}),
    .f({_al_u3105_o,_al_u3103_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u3106|_al_u3097  (
    .a({_al_u3097_o,open_n21254}),
    .b({_al_u3100_o,_al_u1783_o}),
    .c({_al_u3102_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u3105_o,_al_u3096_o}),
    .f({_al_u3106_o,_al_u3097_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B*~A))"),
    //.LUT1("(A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b1111111000000000),
    .INIT_LUT1(16'b1111111011101000),
    .MODE("LOGIC"))
    \_al_u3107|_al_u3424  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 }),
    .f({_al_u3107_o,_al_u3424_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D))"),
    //.LUTF1("(~B*(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D))"),
    //.LUTG0("(B*(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D))"),
    //.LUTG1("(~B*(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D))"),
    .INIT_LUTF0(16'b0000100010001100),
    .INIT_LUTF1(16'b0000001000100011),
    .INIT_LUTG0(16'b0000100010001100),
    .INIT_LUTG1(16'b0000001000100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3108|_al_u3109  (
    .a({_al_u916_o,_al_u1383_o}),
    .b({_al_u3107_o,_al_u3108_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 }),
    .f({_al_u3108_o,_al_u3109_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(~C*B*A))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111111100001000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3111|_al_u3112  (
    .a({open_n21319,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 }),
    .b({open_n21320,_al_u3106_o}),
    .c({_al_u3110_o,_al_u3111_o}),
    .d({_al_u3109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({_al_u3111_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3113|_al_u3110  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u3110_o,_al_u609_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ,_al_u3110_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~C*B))"),
    //.LUT1("(~B*~(~D*~C*A))"),
    .INIT_LUT0(16'b1010001010101010),
    .INIT_LUT1(16'b0011001100110001),
    .MODE("LOGIC"))
    \_al_u3114|_al_u3116  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwuow6_lutinv ,_al_u3114_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ,_al_u3115_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3114_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*~A)))"),
    //.LUT1("(C*~B*D)"),
    .INIT_LUT0(16'b0000000100001111),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"))
    \_al_u3115|_al_u6837  (
    .a({open_n21385,_al_u1269_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,_al_u2868_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u2868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3115_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~B*~(C*A)))"),
    //.LUTF1("(~A*~(D*~(~C*~B)))"),
    //.LUTG0("(D*~(~B*~(C*A)))"),
    //.LUTG1("(~A*~(D*~(~C*~B)))"),
    .INIT_LUTF0(16'b1110110000000000),
    .INIT_LUTF1(16'b0000000101010101),
    .INIT_LUTG0(16'b1110110000000000),
    .INIT_LUTG1(16'b0000000101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3117|_al_u4017  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iugiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .b({_al_u932_o,_al_u903_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .d({_al_u2813_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv }),
    .f({_al_u3117_o,_al_u4017_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u3118|_al_u607  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u3118_o,_al_u607_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(A)*~(D)+(C*B)*A*~(D)+~((C*B))*A*D+(C*B)*A*D)"),
    //.LUTF1("(A*~(D*~(C*~B)))"),
    //.LUTG0("~((C*B)*~(A)*~(D)+(C*B)*A*~(D)+~((C*B))*A*D+(C*B)*A*D)"),
    //.LUTG1("(A*~(D*~(C*~B)))"),
    .INIT_LUTF0(16'b0101010100111111),
    .INIT_LUTF1(16'b0010000010101010),
    .INIT_LUTG0(16'b0101010100111111),
    .INIT_LUTG1(16'b0010000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3120|_al_u3119  (
    .a({_al_u3117_o,_al_u679_o}),
    .b({_al_u3118_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({_al_u3119_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3120_o,_al_u3119_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*~C*B))"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .INIT_LUT0(16'b1010101010100010),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"))
    \_al_u3125|_al_u3126  (
    .a({_al_u1803_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ,_al_u679_o}),
    .c({_al_u3124_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0vow6 ,_al_u3126_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(D*C*~(~B*~A))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b1110000000000000),
    .MODE("LOGIC"))
    \_al_u3129|_al_u3799  (
    .a({_al_u604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u3129_o,_al_u3799_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(~D*~C*B*A)"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"))
    \_al_u3130|_al_u3127  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv }),
    .b({_al_u3126_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u3127_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u3129_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ,_al_u3127_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*B)*~(~D*A))"),
    //.LUT1("(C*A*~(D*~B))"),
    .INIT_LUT0(16'b1111001101010001),
    .INIT_LUT1(16'b1000000010100000),
    .MODE("LOGIC"))
    \_al_u3132|_al_u3131  (
    .a({_al_u3121_o,_al_u1887_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3132_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*C*~A))"),
    //.LUTF1("(~A*(~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    //.LUTG0("(~B*~(D*C*~A))"),
    //.LUTG1("(~A*(~(B)*C*~(D)+B*~(C)*D+~(B)*C*D))"),
    .INIT_LUTF0(16'b0010001100110011),
    .INIT_LUTF1(16'b0001010000010000),
    .INIT_LUTG0(16'b0010001100110011),
    .INIT_LUTG1(16'b0001010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3133|_al_u3134  (
    .a({_al_u1906_o,_al_u3132_o}),
    .b({_al_u1299_o,_al_u3133_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u3133_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("~(~C*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"))
    \_al_u3135|_al_u5009  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 ,\u_cmsdk_mcu/HTRANS [1]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n590 ,_al_u5009_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3136|_al_u404  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3146|_al_u915  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ,_al_u914_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u3147|_al_u3096  (
    .b({open_n21654,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ,_al_u3096_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u3148|_al_u2852  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ,open_n21675}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv ,open_n21676}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Glaiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .d({_al_u1342_o,_al_u1342_o}),
    .f({_al_u3148_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3149|_al_u3192  (
    .b({_al_u1781_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,_al_u606_o}),
    .f({_al_u3149_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~A*~(D*B)))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(C*~(~A*~(D*B)))"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b1110000010100000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1110000010100000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3152|_al_u3151  (
    .a({_al_u3148_o,_al_u609_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yavow6 ,_al_u3150_o}),
    .c({_al_u3149_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u3151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u3152_o,_al_u3151_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3153|_al_u3644  (
    .c({_al_u1346_o,_al_u903_o}),
    .d({_al_u3109_o,_al_u3109_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(~C*~(D*~(~B*~A)))"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(~C*~(D*~(~B*~A)))"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0000000100001111),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0000000100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3154|_al_u4053  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv ,open_n21771}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ,_al_u903_o}),
    .c({_al_u1264_o,_al_u1264_o}),
    .d({_al_u1266_o,_al_u4049_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3156|_al_u3155  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ,open_n21798}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u1269_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }),
    .f({_al_u3156_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3159|_al_u1803  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,open_n21821}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u1803_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u3159_o,_al_u1803_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(~D*C))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001000100000001),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3161|_al_u3160  (
    .a({open_n21842,_al_u3157_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 ,_al_u3158_o}),
    .c({_al_u3160_o,_al_u3159_o}),
    .d({_al_u3152_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ,_al_u3160_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3165|_al_u3164  (
    .a({open_n21863,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F1jiu6_lutinv ,_al_u909_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .d({_al_u3164_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u3165_o,_al_u3164_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~D*C*B))"),
    //.LUT1("(C*A*~(D*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0010000010100000),
    .MODE("LOGIC"))
    \_al_u3167|_al_u3166  (
    .a({_al_u3165_o,_al_u904_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ,_al_u609_o}),
    .c({_al_u3166_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u3167_o,_al_u3166_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3168|_al_u1645  (
    .c({_al_u903_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .d({_al_u609_o,_al_u903_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(D*C))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*~A*~(D*C))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000100010001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000100010001),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3169|_al_u3563  (
    .a({open_n21928,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 }),
    .b({open_n21929,_al_u3186_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u3169_o,_al_u3563_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3170|_al_u3754  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }),
    .f({_al_u3170_o,_al_u3754_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3172|_al_u3171  (
    .a({_al_u3169_o,open_n21982}),
    .b({_al_u3170_o,open_n21983}),
    .c({_al_u1806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~B*A)"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(D*C*~B*A)"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3174|_al_u3173  (
    .a({_al_u3167_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1jiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u3173_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u3174_o,_al_u3173_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~A*~(~C*~B))"),
    //.LUTF1("(D*~(~B*~(C*A)))"),
    //.LUTG0("(D*~A*~(~C*~B))"),
    //.LUTG1("(D*~(~B*~(C*A)))"),
    .INIT_LUTF0(16'b0101010000000000),
    .INIT_LUTF1(16'b1110110000000000),
    .INIT_LUTG0(16'b0101010000000000),
    .INIT_LUTG1(16'b1110110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3176|_al_u3175  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ,_al_u1812_o}),
    .b({_al_u3175_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 }),
    .c({_al_u2373_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3176_o,_al_u3175_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~(B@A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~C*~(B@A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001001),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3178|_al_u6312  (
    .a({open_n22056,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 }),
    .b({open_n22057,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ,_al_u6312_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(~B*~(~D*~C*A))"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(~B*~(~D*~C*A))"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0011001100110001),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0011001100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3180|_al_u3179  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ,open_n22082}),
    .b({_al_u3176_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .c({_al_u3179_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 }),
    .f({_al_u3180_o,_al_u3179_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(A*~(D*B)))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000110100000101),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u3181|_al_u3182  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1jiu6 ,_al_u3181_o}),
    .b({_al_u3174_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0jiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u3180_o,_al_u678_o}),
    .f({_al_u3181_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u3183|_al_u2361  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .d({_al_u2361_o,_al_u1812_o}),
    .f({_al_u3183_o,_al_u2361_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3185|_al_u3184  (
    .b({open_n22153,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv }),
    .c({_al_u3184_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({_al_u3183_o,_al_u1269_o}),
    .f({_al_u3185_o,_al_u3184_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3186|_al_u4153  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv }),
    .c({_al_u1813_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u1812_o,_al_u1813_o}),
    .f({_al_u3186_o,_al_u4153_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3187|_al_u4161  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ,_al_u1582_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .f({_al_u3187_o,_al_u4161_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~(~C*~B)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(A*~(~D*~(~C*~B)))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1010101000000010),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3189|_al_u3627  (
    .a({open_n22228,_al_u3626_o}),
    .b({open_n22229,_al_u3110_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,_al_u903_o}),
    .d({_al_u3110_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u3189_o,_al_u3627_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u3190|_al_u3188  (
    .b({_al_u3189_o,_al_u3187_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 ,_al_u3186_o}),
    .f({_al_u3190_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3191|_al_u3158  (
    .b({open_n22278,_al_u606_o}),
    .c({_al_u696_o,_al_u2829_o}),
    .d({_al_u681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .f({_al_u3191_o,_al_u3158_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(~(D*B)*~(~C*A))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(~(D*B)*~(~C*A))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b0011000111110101),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b0011000111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3194|_al_u3193  (
    .a({_al_u3191_o,_al_u604_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 ,_al_u1907_o}),
    .c({_al_u3193_o,_al_u2392_o}),
    .d({_al_u1582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx9ow6 ,_al_u3193_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(~D*~A)))"),
    //.LUTF1("(C*B*~(D*A))"),
    //.LUTG0("(C*~(B*~(~D*~A)))"),
    //.LUTG1("(C*B*~(D*A))"),
    .INIT_LUTF0(16'b0011000001110000),
    .INIT_LUTF1(16'b0100000011000000),
    .INIT_LUTG0(16'b0011000001110000),
    .INIT_LUTG1(16'b0100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3196|_al_u3195  (
    .a({_al_u3185_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .b({_al_u3190_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx9ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv9ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u3196_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv9ow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3198|_al_u3197  (
    .a({open_n22347,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({_al_u3197_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u3198_o,_al_u3197_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u3200|_al_u3177  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,open_n22370}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3201|_al_u4159  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 ,open_n22391}),
    .b({_al_u679_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbbow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv }),
    .f({_al_u3201_o,_al_u4159_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~B*A*~(D*C))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"))
    \_al_u3203|_al_u3202  (
    .a({_al_u3196_o,open_n22416}),
    .b({_al_u3199_o,open_n22417}),
    .c({_al_u3202_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,_al_u3201_o}),
    .f({_al_u3203_o,_al_u3202_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3205|_al_u2383  (
    .b({_al_u3184_o,open_n22440}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ,_al_u1812_o}),
    .f({_al_u3205_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3206|_al_u3204  (
    .b({_al_u3205_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({_al_u2767_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 ,_al_u1801_o}),
    .f({_al_u3206_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(B*A*~(D*~C))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1000000010001000),
    .MODE("LOGIC"))
    \_al_u3208|_al_u4320  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ,open_n22487}),
    .b({_al_u2771_o,_al_u2365_o}),
    .c({_al_u2370_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 }),
    .f({_al_u3208_o,_al_u4320_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"))
    \_al_u3209|_al_u2754  (
    .a({_al_u2754_o,open_n22508}),
    .b({_al_u1818_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u3149_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 ,_al_u2754_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*A*~(~D*B))"),
    //.LUT1("(D*~C*B*A)"),
    .INIT_LUT0(16'b0000101000000010),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"))
    \_al_u3210|_al_u3613  (
    .a({_al_u3203_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 }),
    .b({_al_u3206_o,_al_u3185_o}),
    .c({_al_u3208_o,_al_u3612_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3210_o,_al_u3613_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3211|_al_u3199  (
    .b({open_n22551,_al_u3198_o}),
    .c({_al_u1269_o,_al_u1269_o}),
    .d({_al_u3183_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 }),
    .f({_al_u3211_o,_al_u3199_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3213|_al_u3212  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u3211_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C*B))"),
    //.LUTF1("(~B*~(A*~(~D*~C)))"),
    //.LUTG0("(A*~(D*~C*B))"),
    //.LUTG1("(~B*~(A*~(~D*~C)))"),
    .INIT_LUTF0(16'b1010001010101010),
    .INIT_LUTF1(16'b0001000100010011),
    .INIT_LUTG0(16'b1010001010101010),
    .INIT_LUTG1(16'b0001000100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3216|_al_u3217  (
    .a({_al_u3214_o,_al_u3216_o}),
    .b({_al_u3215_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({_al_u3216_o,_al_u3217_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~C*B))"),
    //.LUTF1("(A*~(D*~C*B))"),
    //.LUTG0("(A*~(~D*~C*B))"),
    //.LUTG1("(A*~(D*~C*B))"),
    .INIT_LUTF0(16'b1010101010100010),
    .INIT_LUTF1(16'b1010001010101010),
    .INIT_LUTG0(16'b1010101010100010),
    .INIT_LUTG1(16'b1010001010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3219|_al_u3218  (
    .a({_al_u3210_o,_al_u3217_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ,_al_u2380_o}),
    .c({_al_u3218_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u3219_o,_al_u3218_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~D*~C*B))"),
    //.LUTF1("(A*~(D*C*B))"),
    //.LUTG0("(~A*~(~D*~C*B))"),
    //.LUTG1("(A*~(D*C*B))"),
    .INIT_LUTF0(16'b0101010101010001),
    .INIT_LUTF1(16'b0010101010101010),
    .INIT_LUTG0(16'b0101010101010001),
    .INIT_LUTG1(16'b0010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3224|_al_u3222  (
    .a({_al_u3222_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hs8ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 }),
    .c({_al_u3223_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u3124_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .f({_al_u3224_o,_al_u3222_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~B*D))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000110000001111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u3226|_al_u3225  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,open_n22670}),
    .b({_al_u912_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({_al_u3225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }),
    .f({_al_u3226_o,_al_u3225_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3227|_al_u2386  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u2364_o,_al_u2364_o}),
    .f({_al_u3227_o,_al_u2386_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~A*~(~C*B)))"),
    //.LUT1("(~A*~(D*C*B))"),
    .INIT_LUT0(16'b0000000010101110),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"))
    \_al_u3229|_al_u3228  (
    .a({_al_u3226_o,_al_u3227_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xz9ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u1269_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xz9ow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*~(D*~A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*~(D*~A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000011000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3230|_al_u3221  (
    .a({_al_u3221_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 }),
    .b({_al_u3224_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv }),
    .c({_al_u3229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u3230_o,_al_u3221_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3231|_al_u3233  (
    .a({open_n22759,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 }),
    .b({open_n22760,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 }),
    .d({_al_u2771_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 ,_al_u3233_o}));
  // ../RTL/cortexm0ds_logic.v(17747)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*C)*~(~B*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110100001101),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3235|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6_reg  (
    .a({_al_u3219_o,_al_u3235_o}),
    .b({_al_u3230_o,_al_u3240_o}),
    .c({_al_u3233_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u3234_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3235_o,open_n22794}),
    .q({open_n22798,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }));  // ../RTL/cortexm0ds_logic.v(17747)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(~D*A))"),
    //.LUTF1("(~(C*B)*~(~D*A))"),
    //.LUTG0("(~(~C*B)*~(~D*A))"),
    //.LUTG1("(~(C*B)*~(~D*A))"),
    .INIT_LUTF0(16'b1111001101010001),
    .INIT_LUTF1(16'b0011111100010101),
    .INIT_LUTG0(16'b1111001101010001),
    .INIT_LUTG1(16'b0011111100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3238|_al_u3237  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 ,_al_u1271_o}),
    .b({_al_u681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 }),
    .c({_al_u3236_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u3237_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3238_o,_al_u3237_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(D*~(A*~(C*B)))"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(D*~(A*~(C*B)))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1101010100000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b1101010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3240|_al_u3239  (
    .a({_al_u3238_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ,_al_u604_o}),
    .c({_al_u3239_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u3109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u3240_o,_al_u3239_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3244|_al_u3854  (
    .b({open_n22849,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({_al_u2763_o,_al_u2763_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ,_al_u3854_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3245|_al_u3307  (
    .b({_al_u2759_o,_al_u2759_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv }),
    .f({_al_u3245_o,_al_u3307_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u3247|_al_u3246  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,open_n22902}),
    .c({_al_u3246_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u912_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ,_al_u3246_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(D*C*~B*A)"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3249|_al_u3242  (
    .a({_al_u3242_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv }),
    .b({_al_u3243_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 }),
    .c({_al_u3245_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({_al_u3248_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .f({_al_u3249_o,_al_u3242_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(A@(D*C)))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~B*(A@(D*C)))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001001000100010),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001000100010),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3250|_al_u2791  (
    .a({open_n22947,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,_al_u2790_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S88iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 ,_al_u2791_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(B@(A*C*~(D)+A*~(C)*D+~(A)*C*D+A*C*D))"),
    .INIT_LUT0(16'b0111111011101000),
    .INIT_LUT1(16'b0011011001101100),
    .MODE("LOGIC"))
    \_al_u3252|_al_u3251  (
    .a({_al_u2785_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17402)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(A*~(D*~C)))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(~B*~(A*~(D*~C)))"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110110011101110),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1110110011101110),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3255|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6_reg  (
    .a({open_n22992,_al_u2467_o}),
    .b({open_n22993,_al_u2468_o}),
    .c({_al_u2468_o,_al_u2469_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U73iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u2467_o,_al_u2470_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u3255_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 }),
    .q({open_n23013,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gylpw6 }));  // ../RTL/cortexm0ds_logic.v(17402)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*~A)"),
    //.LUTF1("(~D*C*B*~A)"),
    //.LUTG0("(~D*C*B*~A)"),
    //.LUTG1("(~D*C*B*~A)"),
    .INIT_LUTF0(16'b0000000001000000),
    .INIT_LUTF1(16'b0000000001000000),
    .INIT_LUTG0(16'b0000000001000000),
    .INIT_LUTG1(16'b0000000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3257|_al_u3776  (
    .a({_al_u3255_o,_al_u3255_o}),
    .b({_al_u3256_o,_al_u1757_o}),
    .c({_al_u1250_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ,_al_u3776_o}));
  // ../RTL/cortexm0ds_logic.v(17383)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3259|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6_reg  (
    .c({_al_u3258_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ,_al_u3259_o}),
    .mi({open_n23045,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .f({_al_u3259_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 }),
    .q({open_n23061,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }));  // ../RTL/cortexm0ds_logic.v(17383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3267|_al_u400  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3270|_al_u519  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] }),
    .f({_al_u3270_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3271|_al_u3335  (
    .c({_al_u1772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv }),
    .d({_al_u3270_o,_al_u3270_o}),
    .f({_al_u3271_o,_al_u3335_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3275|_al_u3287  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 }),
    .f({_al_u3275_o,_al_u3287_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3276|_al_u3734  (
    .a({open_n23158,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv }),
    .b({open_n23159,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 }),
    .d({_al_u3275_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ,_al_u3734_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3280|_al_u1772  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] }),
    .f({_al_u3280_o,_al_u1772_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3281|_al_u3372  (
    .c({_al_u3280_o,_al_u1772_o}),
    .d({_al_u3275_o,_al_u3275_o}),
    .f({_al_u3281_o,_al_u3372_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3288|_al_u3436  (
    .c({_al_u3280_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv }),
    .d({_al_u3287_o,_al_u3287_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~A*(C@(D*B)))"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~A*(C@(D*B)))"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0001010001010000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0001010001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3306|_al_u6042  (
    .a({_al_u2783_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .f({_al_u3306_o,_al_u6042_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3308|_al_u1371  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ,open_n23284}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ,open_n23285}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .f({_al_u3308_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D*~A))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(~(C*~B)*~(D*~A))"),
    //.LUTG1("(D*C*~B*A)"),
    .INIT_LUTF0(16'b1000101011001111),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b1000101011001111),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3309|_al_u3305  (
    .a({_al_u3305_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hd8iu6_lutinv }),
    .b({_al_u3306_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 }),
    .c({_al_u3307_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .d({_al_u3308_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({_al_u3309_o,_al_u3305_o}));
  // ../RTL/cortexm0ds_logic.v(17419)
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(~C*(D@B)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(A*~(~C*(D@B)))"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101011101011101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0101011101011101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3310|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6_reg  (
    .a({open_n23334,_al_u3249_o}),
    .b({open_n23335,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv ,_al_u2790_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7biu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 ,open_n23353}),
    .q({open_n23357,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 }));  // ../RTL/cortexm0ds_logic.v(17419)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u3313|_al_u3312  (
    .a({open_n23358,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .d({_al_u3312_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({_al_u3313_o,_al_u3312_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B@(A*C*~(D)+A*~(C)*D+~(A)*C*D+A*C*D))"),
    //.LUT1("(A*~(D*C*B))"),
    .INIT_LUT0(16'b0011011001101100),
    .INIT_LUT1(16'b0010101010101010),
    .MODE("LOGIC"))
    \_al_u3314|_al_u3253  (
    .a({_al_u3313_o,_al_u2786_o}),
    .b({_al_u2786_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3314_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7biu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    .INIT_LUT0(16'b1111000000001111),
    .MODE("LOGIC"))
    _al_u3315 (
    .c({open_n23403,_al_u3314_o}),
    .d({open_n23406,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv }),
    .f({open_n23420,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gcjiu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A*~(C@B))"),
    //.LUT1("(~D*(C@B))"),
    .INIT_LUT0(16'b0000000001000001),
    .INIT_LUT1(16'b0000000000111100),
    .MODE("LOGIC"))
    \_al_u3317|_al_u3258  (
    .a({open_n23426,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv ,_al_u3258_o}));
  // ../RTL/cortexm0ds_logic.v(18013)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(D*C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3318|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 ,open_n23447}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi1iu6_lutinv }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 ,_al_u3872_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u3318_o,open_n23465}),
    .q({open_n23469,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ry2qw6 }));  // ../RTL/cortexm0ds_logic.v(18013)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3320|_al_u3882  (
    .b({open_n23472,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph1iu6 }),
    .c({_al_u3319_o,_al_u3319_o}),
    .d({_al_u3318_o,_al_u3318_o}),
    .f({_al_u3320_o,_al_u3882_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u3322|_al_u3869  (
    .a({_al_u3255_o,open_n23493}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv ,_al_u3255_o}),
    .f({_al_u3322_o,_al_u3869_o}));
  // ../RTL/cortexm0ds_logic.v(17597)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~(D*~(A)*~((C*B))+D*A*~((C*B))+~(D)*A*(C*B)+D*A*(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100000001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3324|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6_reg  (
    .a({\u_cmsdk_mcu/dbg_swdo ,open_n23514}),
    .b({_al_u1676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 }),
    .mi({open_n23525,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 }),
    .f({_al_u3324_o,\u_cmsdk_mcu/dbg_swdo }),
    .q({open_n23530,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 }));  // ../RTL/cortexm0ds_logic.v(17597)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~C*~B*~D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3327|_al_u3326  (
    .b({_al_u3326_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .c({_al_u1757_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ,_al_u529_o}),
    .f({_al_u3327_o,_al_u3326_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(D*~B*~(~C*A))"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0011000100000000),
    .MODE("LOGIC"))
    \_al_u3329|_al_u1759  (
    .a({_al_u3327_o,open_n23557}),
    .b({_al_u530_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .c({_al_u3328_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ,_al_u1758_o}),
    .f({_al_u3329_o,_al_u1759_o}));
  // ../RTL/cortexm0ds_logic.v(17333)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(D)*~(B)*~(C)+~(D)*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(D)*~(B)*~(C)+~(D)*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b1111000011001111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b1111000011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3330|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6_reg  (
    .b({_al_u3329_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/It3iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u3325_o,_al_u3323_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/It3iu6_lutinv ,open_n23598}),
    .q({open_n23602,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 }));  // ../RTL/cortexm0ds_logic.v(17333)
  // ../RTL/cortexm0ds_logic.v(17598)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~(C*B)))"),
    //.LUT1("(~(~D*C)*~(B*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000010101010),
    .INIT_LUT1(16'b0111011100000111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3333|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6_reg  (
    .a({\u_cmsdk_mcu/HWDATA [0],_al_u3333_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ,\u_cmsdk_mcu/HWDATA [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 }),
    .mi({open_n23613,\u_cmsdk_mcu/HWDATA [0]}),
    .f({_al_u3333_o,_al_u3334_o}),
    .q({open_n23618,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 }));  // ../RTL/cortexm0ds_logic.v(17598)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(D*~A))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1000000011000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3337|_al_u480  (
    .a({open_n23619,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_overrun ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .f({_al_u3337_o,_al_u480_o}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~(C*B)))"),
    //.LUT1("(~(~D*~C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000010101010),
    .INIT_LUT1(16'b0111011101110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3338|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b8  (
    .a({\u_cmsdk_mcu/HWDATA [8],_al_u3338_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ,\u_cmsdk_mcu/HWDATA [8]}),
    .c({_al_u3337_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 }),
    .mi({open_n23650,\u_cmsdk_mcu/HWDATA [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3338_o,_al_u3339_o}),
    .q({open_n23654,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [8]}));  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3343|_al_u3362  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv }),
    .d({_al_u3270_o,_al_u3275_o}),
    .f({_al_u3343_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3346|_al_u3340  (
    .c({_al_u1772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv }),
    .d({_al_u3287_o,_al_u3287_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3350|_al_u3446  (
    .b({_al_u3280_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ,_al_u1772_o}),
    .f({_al_u3350_o,_al_u3446_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3353|_al_u3443  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ,_al_u3443_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3355|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12],open_n23755}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [14]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [14]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n299 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3355_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [14]}),
    .q({open_n23771,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u3356|_al_u3952  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0],open_n23772}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1],_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv }),
    .f({_al_u3356_o,_al_u3952_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3357|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6],open_n23793}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n285 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3357_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [7]}),
    .q({open_n23809,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3358|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2],open_n23810}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [5]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n281 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3358_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [5]}),
    .q({open_n23830,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3359|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b6  (
    .a({_al_u3355_o,open_n23831}),
    .b({_al_u3356_o,open_n23832}),
    .c({_al_u3357_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6]}),
    .clk(1'b1),
    .d({_al_u3358_o,_al_u3068_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3359_o,open_n23846}),
    .q({open_n23850,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [6]}));  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u3365|_al_u4876  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [13]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[13] }),
    .f({_al_u3365_o,_al_u4876_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3366|_al_u3534  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] ,open_n23871}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [6]}),
    .f({_al_u3366_o,_al_u3534_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3367|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] ,open_n23896}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] ,open_n23897}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n285 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3367_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [7]}),
    .q({open_n23913,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3368|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] ,open_n23914}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] ,open_n23915}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n281 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3368_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [5]}),
    .q({open_n23935,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3369|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b7  (
    .a({_al_u3365_o,open_n23936}),
    .b({_al_u3366_o,open_n23937}),
    .c({_al_u3367_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7]}),
    .clk(1'b1),
    .d({_al_u3368_o,_al_u3073_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3369_o,open_n23955}),
    .q({open_n23959,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [7]}));  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3374|_al_u521  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3377|_al_u3376  (
    .b({open_n23988,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] }),
    .c({_al_u1772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 }));
  // ../RTL/cortexm0ds_logic.v(17682)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(C*~(D*~B)))"),
    //.LUT1("(C*~(B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101010111110101),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3378|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6_reg  (
    .a({open_n24013,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ,_al_u2721_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ,_al_u3378_o}),
    .clk(XTAL1_wire),
    .d({_al_u1777_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3378_o,open_n24027}),
    .q({open_n24031,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 }));  // ../RTL/cortexm0ds_logic.v(17682)
  // ../RTL/cortexm0ds_logic.v(17435)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTG1("(C*~(B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011001111110000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1011001111110000),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3381|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6_reg  (
    .a({open_n24032,_al_u2729_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ,_al_u2733_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ,_al_u3381_o}),
    .clk(XTAL1_wire),
    .d({_al_u1777_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3381_o,open_n24050}),
    .q({open_n24054,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 }));  // ../RTL/cortexm0ds_logic.v(17435)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*~D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"))
    \_al_u3385|_al_u3384  (
    .a({open_n24055,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv ,_al_u2299_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .d({_al_u3384_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 }),
    .f({_al_u3385_o,_al_u3384_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u3387|_al_u2296  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({_al_u2296_o,_al_u1251_o}),
    .f({_al_u3387_o,_al_u2296_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3390|_al_u3389  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .d({_al_u529_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epyhu6 }),
    .f({_al_u3390_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A*~(C*B))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~D*~A*~(C*B))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000000000010101),
    .INIT_LUTF1(16'b1111010100010011),
    .INIT_LUTG0(16'b0000000000010101),
    .INIT_LUTG1(16'b1111010100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3391|_al_u4272  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ,_al_u2299_o}),
    .b({_al_u3390_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .f({_al_u3391_o,_al_u4272_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C*B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~(D*C*B))"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b0010101010101010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0010101010101010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3392|_al_u3388  (
    .a({_al_u3388_o,_al_u3387_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ,_al_u1308_o}),
    .c({_al_u3391_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .d({_al_u2305_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .f({_al_u3392_o,_al_u3388_o}));
  // ../RTL/cortexm0ds_logic.v(17338)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D*~(B*~A)))"),
    //.LUT1("(~D*(C@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101111110000),
    .INIT_LUT1(16'b0000000000111100),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3393|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6_reg  (
    .a({open_n24168,_al_u3385_o}),
    .b({_al_u529_o,_al_u3392_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 ,_al_u3393_o}),
    .clk(SWCLKTCK_pad),
    .d({_al_u1761_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u3393_o,open_n24182}),
    .q({open_n24186,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }));  // ../RTL/cortexm0ds_logic.v(17338)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3396|_al_u3395  (
    .b({_al_u3395_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }),
    .c({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u1775_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u3396_o,_al_u3395_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(A*~(D*B)))"),
    //.LUTF1("(B*A*~(~D*C))"),
    //.LUTG0("(~C*~(A*~(D*B)))"),
    //.LUTG1("(B*A*~(~D*C))"),
    .INIT_LUTF0(16'b0000110100000101),
    .INIT_LUTF1(16'b1000100000001000),
    .INIT_LUTG0(16'b0000110100000101),
    .INIT_LUTG1(16'b1000100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3398|_al_u3399  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epjiu6 ,_al_u3398_o}),
    .b({_al_u3397_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hviiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,_al_u609_o}),
    .f({_al_u3398_o,_al_u3399_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~C*~B*~(D*A))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000000100000011),
    .MODE("LOGIC"))
    \_al_u3400|_al_u2836  (
    .a({_al_u2771_o,_al_u2365_o}),
    .b({_al_u2773_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({_al_u2836_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({_al_u3400_o,_al_u2836_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(A*~(~C*~(~D*~B)))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(A*~(~C*~(~D*~B)))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1010000010100010),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1010000010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3402|_al_u3401  (
    .a({_al_u3400_o,open_n24257}),
    .b({_al_u3401_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u909_o,_al_u2365_o}),
    .f({_al_u3402_o,_al_u3401_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u3403|_al_u3410  (
    .a({open_n24282,_al_u3402_o}),
    .b({open_n24283,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 }),
    .c({_al_u2771_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({_al_u3402_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ,_al_u3410_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3404|_al_u4410  (
    .b({_al_u912_o,_al_u2832_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({_al_u2832_o,_al_u2771_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ,_al_u4410_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"))
    \_al_u3405|_al_u3554  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ,open_n24326}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .f({_al_u3405_o,_al_u3554_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3406|_al_u3558  (
    .b({open_n24349,_al_u604_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dr7ow6 ,_al_u3558_o}));
  // ../RTL/cortexm0ds_logic.v(18705)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUTG1("(C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011111110010),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b1111011111110010),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3408|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6_reg  (
    .a({open_n24374,_al_u3399_o}),
    .b({_al_u1383_o,_al_u3405_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6iow6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6iow6_lutinv ,open_n24393}),
    .q({open_n24397,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umkax6 }));  // ../RTL/cortexm0ds_logic.v(18705)
  // ../RTL/cortexm0ds_logic.v(18634)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUT1("(C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011111110010),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3411|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6_reg  (
    .a({open_n24398,_al_u3399_o}),
    .b({_al_u1765_o,_al_u3410_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkhow6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkhow6_lutinv ,open_n24413}),
    .q({open_n24417,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6jax6 }));  // ../RTL/cortexm0ds_logic.v(18634)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*~(~C*~B*~A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*~(~C*~B*~A))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111111000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111111000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3413|_al_u906  (
    .a({_al_u906_o,open_n24418}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ,open_n24419}),
    .c({_al_u1359_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 ,_al_u906_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u3415|_al_u3414  (
    .a({open_n24444,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 }),
    .d({_al_u3414_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u3415_o,_al_u3414_o}));
  // ../RTL/cortexm0ds_logic.v(17625)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011111110010),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3417|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ,_al_u3399_o}),
    .b({_al_u916_o,_al_u3416_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pj7ow6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pj7ow6_lutinv ,open_n24479}),
    .q({open_n24483,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fkrpw6 }));  // ../RTL/cortexm0ds_logic.v(17625)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u3420|_al_u3419  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmiiu6 ,open_n24484}),
    .b({_al_u2832_o,open_n24485}),
    .c({_al_u3419_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({_al_u3420_o,_al_u3419_o}));
  // ../RTL/cortexm0ds_logic.v(18704)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUT1("(D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011111110010),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3422|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6_reg  (
    .a({open_n24506,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljiiu6 ,_al_u3422_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoiiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({_al_u3421_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 }),
    .f({_al_u3422_o,open_n24521}),
    .q({open_n24525,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 }));  // ../RTL/cortexm0ds_logic.v(18704)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3425|_al_u3423  (
    .b({open_n24528,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({_al_u3424_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u3423_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoiiu6_lutinv ,_al_u3423_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~C*B*~(D*~A))"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0000100000001100),
    .MODE("LOGIC"))
    \_al_u3429|_al_u3328  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv ,_al_u1251_o}),
    .b({_al_u3391_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .c({_al_u3328_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .f({_al_u3429_o,_al_u3328_o}));
  // ../RTL/cortexm0ds_logic.v(17374)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(~D*C*~A))"),
    //.LUT1("(B*~(C*~D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001101110011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3431|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6_reg  (
    .a({open_n24573,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmyhu6 }),
    .b({_al_u3430_o,_al_u3431_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ,_al_u1253_o}),
    .clk(SWCLKTCK_pad),
    .d({_al_u3429_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u3431_o,open_n24587}),
    .q({open_n24591,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }));  // ../RTL/cortexm0ds_logic.v(17374)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~A*~(C*B)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~D*~(~A*~(C*B)))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000011101010),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000011101010),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3433|_al_u1024  (
    .a({open_n24592,_al_u1020_o}),
    .b({open_n24593,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [0],_al_u1023_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [10],_al_u1024_o}));
  // ../RTL/cortexm0ds_logic.v(19299)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0101111100010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3434|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6_reg  (
    .a({\u_cmsdk_mcu/HWDATA [10],open_n24618}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [10],open_n24619}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ,_al_u3938_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3434_o,open_n24633}),
    .q({open_n24637,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 }));  // ../RTL/cortexm0ds_logic.v(19299)
  // ../RTL/cortexm0ds_logic.v(19305)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(A*~(D*~(C*B)))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(A*~(D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1000000010101010),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3435|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6_reg  (
    .a({_al_u3434_o,open_n24638}),
    .b({\u_cmsdk_mcu/HWDATA [10],_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ,_al_u3435_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3435_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3phu6 }),
    .q({open_n24659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 }));  // ../RTL/cortexm0ds_logic.v(19305)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3438|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [4],open_n24660}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [2],open_n24661}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2],_al_u2496_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4],\u_cmsdk_mcu/HWDATA [4]}),
    .mi({open_n24672,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3438_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n62 }),
    .q({open_n24676,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4]}));  // ../RTL/gpio_apbif.v(323)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3439|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [5],open_n24677}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [3],open_n24678}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [3],_al_u2496_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5],\u_cmsdk_mcu/HWDATA [3]}),
    .mi({open_n24689,\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3439_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n60 }),
    .q({open_n24693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [3]}));  // ../RTL/gpio_apbif.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3440|_al_u3703  (
    .a({open_n24694,_al_u3699_o}),
    .b({open_n24695,_al_u3700_o}),
    .c({_al_u3439_o,_al_u3701_o}),
    .d({_al_u3438_o,_al_u3702_o}),
    .f({_al_u3440_o,_al_u3703_o}));
  // ../RTL/cortexm0ds_logic.v(19287)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*~B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0101111101001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3441|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6_reg  (
    .a({\u_cmsdk_mcu/HWDATA [12],open_n24716}),
    .b({_al_u3440_o,open_n24717}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ,_al_u3941_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3441_o,open_n24731}),
    .q({open_n24735,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 }));  // ../RTL/cortexm0ds_logic.v(19287)
  // ../RTL/cortexm0ds_logic.v(19293)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(A*~(D*~(C*B)))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(A*~(D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1000000010101010),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3442|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6_reg  (
    .a({_al_u3441_o,open_n24736}),
    .b({\u_cmsdk_mcu/HWDATA [12],_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ,_al_u3443_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ,_al_u3442_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3442_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2phu6 }),
    .q({open_n24757,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 }));  // ../RTL/cortexm0ds_logic.v(19293)
  // ../RTL/cortexm0ds_logic.v(17636)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0010000001110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3445|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6_reg  (
    .a({\u_cmsdk_mcu/HWDATA [15],open_n24758}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ,_al_u3446_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ,_al_u3445_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3445_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1phu6 }),
    .q({open_n24775,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 }));  // ../RTL/cortexm0ds_logic.v(17636)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3450|_al_u635  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1],open_n24778}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]}),
    .f({_al_u3450_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt2/o_1_lutinv }));
  // ../RTL/cortexm0ds_logic.v(19353)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~B*~A*~(~D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0001000100010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3451|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6_reg  (
    .a({_al_u3448_o,open_n24803}),
    .b({_al_u3449_o,_al_u1777_o}),
    .c({_al_u3450_o,_al_u3454_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 ,_al_u3451_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3451_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1phu6 }),
    .q({open_n24820,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 }));  // ../RTL/cortexm0ds_logic.v(19353)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u3452|_al_u3269  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3453|_al_u3463  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ,_al_u3453_o}),
    .f({_al_u3453_o,_al_u3463_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3454|_al_u3468  (
    .c({_al_u3280_o,_al_u1772_o}),
    .d({_al_u3453_o,_al_u3453_o}),
    .f({_al_u3454_o,_al_u3468_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3458|_al_u3931  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 ,_al_u3925_o}),
    .c({_al_u3280_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ,_al_u3931_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(C*~(B*D))"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"))
    \_al_u3460|_al_u3532  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 }),
    .d({\u_cmsdk_mcu/HWDATA [18],\u_cmsdk_mcu/HWDATA [16]}),
    .f({_al_u3460_o,_al_u3532_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3462|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b2  (
    .a({_al_u3460_o,open_n24949}),
    .b({_al_u3461_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [2]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n275 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3462_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [2]}),
    .q({open_n24969,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3467|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b19  (
    .a({_al_u3465_o,open_n24970}),
    .b({_al_u3466_o,open_n24971}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 ,\u_cmsdk_mcu/HWDATA [19]}),
    .mi({open_n24975,\u_cmsdk_mcu/HWDATA [19]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3467_o,_al_u3466_o}),
    .q({open_n24990,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [19]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cortexm0ds_logic.v(19413)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3472|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6_reg  (
    .a({_al_u3470_o,open_n24991}),
    .b({_al_u3471_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 ,_al_u3472_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3472_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0phu6 }),
    .q({open_n25012,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 }));  // ../RTL/cortexm0ds_logic.v(19413)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3473|_al_u3494  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv }),
    .f({_al_u3473_o,_al_u3494_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3474|_al_u3489  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ,_al_u1772_o}),
    .d({_al_u3473_o,_al_u3473_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ,_al_u3489_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3478|_al_u3477  (
    .a({_al_u3476_o,open_n25059}),
    .b({_al_u3477_o,open_n25060}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 ,\u_cmsdk_mcu/HWDATA [21]}),
    .f({_al_u3478_o,_al_u3477_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3479|_al_u3484  (
    .c({_al_u3280_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv }),
    .d({_al_u3473_o,_al_u3473_o}),
    .f({_al_u3479_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(20051)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3483|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6_reg  (
    .a({_al_u3481_o,open_n25109}),
    .b({_al_u3482_o,open_n25110}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 ,\u_cmsdk_mcu/HWDATA [22]}),
    .mi({open_n25114,\u_cmsdk_mcu/HWDATA [22]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3483_o,_al_u3482_o}),
    .q({open_n25129,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 }));  // ../RTL/cortexm0ds_logic.v(20051)
  // ../RTL/cortexm0ds_logic.v(18958)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3488|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6_reg  (
    .a({_al_u3486_o,open_n25130}),
    .b({_al_u3487_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 ,\u_cmsdk_mcu/HWDATA [23]}),
    .mi({open_n25134,\u_cmsdk_mcu/HWDATA [23]}),
    .f({_al_u3488_o,_al_u3486_o}),
    .q({open_n25150,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 }));  // ../RTL/cortexm0ds_logic.v(18958)
  // ../RTL/cortexm0ds_logic.v(19461)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3493|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6_reg  (
    .a({_al_u3491_o,open_n25151}),
    .b({_al_u3492_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 ,_al_u3493_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3493_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdpw6 }),
    .q({open_n25168,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 }));  // ../RTL/cortexm0ds_logic.v(19461)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3495|_al_u3943  (
    .b({open_n25171,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]}),
    .d({_al_u3494_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ,_al_u3943_o}));
  // ../RTL/cortexm0ds_logic.v(19437)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3499|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6_reg  (
    .a({_al_u3497_o,open_n25196}),
    .b({_al_u3498_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 ,_al_u3499_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3499_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwdpw6 }),
    .q({open_n25213,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 }));  // ../RTL/cortexm0ds_logic.v(19437)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3500|_al_u3510  (
    .c({_al_u3280_o,_al_u1772_o}),
    .d({_al_u3494_o,_al_u3494_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(19473)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3504|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6_reg  (
    .a({_al_u3502_o,open_n25242}),
    .b({_al_u3503_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 ,_al_u3504_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzohu6 }),
    .q({open_n25263,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 }));  // ../RTL/cortexm0ds_logic.v(19473)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3505|_al_u3949  (
    .b({open_n25266,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]}),
    .d({_al_u3494_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ,_al_u3949_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3509|_al_u3508  (
    .a({_al_u3507_o,open_n25287}),
    .b({_al_u3508_o,open_n25288}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 ,_al_u2729_o}),
    .f({_al_u3509_o,_al_u3508_o}));
  // ../RTL/cortexm0ds_logic.v(19497)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3514|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6_reg  (
    .a({_al_u3512_o,open_n25313}),
    .b({_al_u3513_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12],_al_u3515_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 ,_al_u3514_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xyohu6 }),
    .q({open_n25330,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 }));  // ../RTL/cortexm0ds_logic.v(19497)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3515|_al_u3955  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ,_al_u3515_o}),
    .f({_al_u3515_o,_al_u3955_o}));
  // ../RTL/cortexm0ds_logic.v(19047)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3519|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6_reg  (
    .a({_al_u3517_o,open_n25357}),
    .b({_al_u3518_o,open_n25358}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 ,\u_cmsdk_mcu/HWDATA [30]}),
    .mi({open_n25369,\u_cmsdk_mcu/HWDATA [30]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3519_o,_al_u3518_o}),
    .q({open_n25373,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 }));  // ../RTL/cortexm0ds_logic.v(19047)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3520|_al_u3525  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv ,_al_u1772_o}),
    .f({_al_u3520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 }));
  // ../RTL/cortexm0ds_logic.v(19593)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3524|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6_reg  (
    .a({_al_u3522_o,open_n25396}),
    .b({_al_u3523_o,open_n25397}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 ,\u_cmsdk_mcu/HWDATA [31]}),
    .mi({open_n25408,\u_cmsdk_mcu/HWDATA [31]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3524_o,_al_u3523_o}),
    .q({open_n25412,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 }));  // ../RTL/cortexm0ds_logic.v(19593)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3529|_al_u3528  (
    .a({_al_u3527_o,open_n25413}),
    .b({_al_u3528_o,open_n25414}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 ,_al_u2741_o}),
    .f({_al_u3529_o,_al_u3528_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3530|_al_u3984  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv ,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]}),
    .d({_al_u3280_o,_al_u3530_o}),
    .f({_al_u3530_o,_al_u3984_o}));
  // ../RTL/cortexm0ds_logic.v(19359)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~A)"),
    //.LUTF1("(~B*~A*~(~D*~C))"),
    //.LUTG0("(D*~C*~B*~A)"),
    //.LUTG1("(~B*~A*~(~D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0001000100010000),
    .INIT_LUTG0(16'b0000000100000000),
    .INIT_LUTG1(16'b0001000100010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3535|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6_reg  (
    .a({_al_u3532_o,_al_u3874_o}),
    .b({_al_u3533_o,_al_u3533_o}),
    .c({_al_u3534_o,_al_u3534_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 ,_al_u3929_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3535_o,open_n25482}),
    .q({open_n25486,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 }));  // ../RTL/cortexm0ds_logic.v(19359)
  EG_PHY_MSLICE #(
    //.LUT0("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011111100001000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3536|_al_u3929  (
    .a({open_n25487,_al_u1777_o}),
    .b({open_n25488,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukbpw6_lutinv ,_al_u3925_o}),
    .d({_al_u3453_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1bx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ,_al_u3929_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B@D))"),
    //.LUTF1("(~D*C*B*~A)"),
    //.LUTG0("(C*~(B@D))"),
    //.LUTG1("(~D*C*B*~A)"),
    .INIT_LUTF0(16'b1100000000110000),
    .INIT_LUTF1(16'b0000000001000000),
    .INIT_LUTG0(16'b1100000000110000),
    .INIT_LUTG1(16'b0000000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3540|_al_u3539  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,open_n25509}),
    .b({_al_u3539_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({_al_u3540_o,_al_u3539_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~A*~(D*~B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"))
    \_al_u3542|_al_u3538  (
    .a({_al_u3538_o,open_n25534}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cn7ow6 ,open_n25535}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtbow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cbbiu6_lutinv }),
    .f({_al_u3542_o,_al_u3538_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C@B@D)"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(C@B@D)"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b1100001100111100),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b1100001100111100),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3543|_al_u2786  (
    .b({_al_u3542_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv ,_al_u2785_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itbow6 ,_al_u2786_o}));
  // ../RTL/cortexm0ds_logic.v(17878)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUTG1("(C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011111110010),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b1111011111110010),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3544|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6_reg  (
    .a({open_n25582,_al_u3399_o}),
    .b({_al_u916_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itbow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,_al_u3544_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk7ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .f({_al_u3544_o,open_n25601}),
    .q({open_n25605,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }));  // ../RTL/cortexm0ds_logic.v(17878)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~(~C*B)))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000100010101010),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u3546|_al_u4390  (
    .a({open_n25606,_al_u4389_o}),
    .b({_al_u2832_o,_al_u2369_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dcziu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eciiu6 ,_al_u4390_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u3548|_al_u3547  (
    .b({_al_u2841_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eciiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({_al_u3547_o,_al_u2827_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbiiu6 ,_al_u3547_o}));
  // ../RTL/cortexm0ds_logic.v(18702)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*(~D*~(B)*~(A)+~D*B*~(A)+~(~D)*B*A+~D*B*A))"),
    //.LUT1("(C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011111110010),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3549|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6_reg  (
    .a({open_n25649,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbiiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ,_al_u3549_o}),
    .clk(XTAL1_wire),
    .d({_al_u3423_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 }),
    .f({_al_u3549_o,open_n25664}),
    .q({open_n25668,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 }));  // ../RTL/cortexm0ds_logic.v(18702)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*~(D*C*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0001001100110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001001100110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3551|_al_u2790  (
    .a({open_n25669,_al_u2771_o}),
    .b({open_n25670,_al_u2789_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yy7ow6 ,_al_u2790_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~A*~(D*C*~B))"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~A*~(D*C*~B))"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0100010101010101),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0100010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3553|_al_u3552  (
    .a({_al_u3552_o,_al_u2771_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yy7ow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({_al_u3553_o,_al_u3552_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(B*~(A*~(D*C)))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1100010001000100),
    .MODE("LOGIC"))
    \_al_u3556|_al_u3555  (
    .a({_al_u3553_o,_al_u2369_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ,_al_u3554_o}),
    .c({_al_u2832_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u3555_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({_al_u3556_o,_al_u3555_o}));
  // ../RTL/cmsdk_apb_uart.v(614)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u355|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b0  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [2],_al_u355_o}),
    .mi({open_n25744,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u355_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc }),
    .q({open_n25759,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [0]}));  // ../RTL/cmsdk_apb_uart.v(614)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~(~D*~A))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~C*B*~(~D*~A))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000110000001000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000110000001000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3561|_al_u3560  (
    .a({_al_u3169_o,_al_u682_o}),
    .b({_al_u3558_o,_al_u1346_o}),
    .c({_al_u3559_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u3560_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3561_o,_al_u3560_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~B*~(~D*C)))"),
    //.LUTF1("(C*A*~(D*B))"),
    //.LUTG0("(A*~(~B*~(~D*C)))"),
    //.LUTG1("(C*A*~(D*B))"),
    .INIT_LUTF0(16'b1000100010101000),
    .INIT_LUTF1(16'b0010000010100000),
    .INIT_LUTG0(16'b1000100010101000),
    .INIT_LUTG1(16'b0010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3564|_al_u3562  (
    .a({_al_u3561_o,_al_u2361_o}),
    .b({_al_u3562_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({_al_u3563_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7kiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u3564_o,_al_u3562_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(A*~(D*B)))"),
    //.LUT1("(D*C*~B*~A)"),
    .INIT_LUT0(16'b1111001011111010),
    .INIT_LUT1(16'b0001000000000000),
    .MODE("LOGIC"))
    \_al_u3565|_al_u3566  (
    .a({_al_u3556_o,_al_u3565_o}),
    .b({_al_u3557_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbiow6_lutinv }),
    .c({_al_u3564_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lv7ow6 ,_al_u678_o}),
    .f({_al_u3565_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u3567|_al_u2408  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~C*A))"),
    //.LUTF1("(~B*A*~(D*C))"),
    //.LUTG0("(~B*~(D*~C*A))"),
    //.LUTG1("(~B*A*~(D*C))"),
    .INIT_LUTF0(16'b0011000100110011),
    .INIT_LUTF1(16'b0000001000100010),
    .INIT_LUTG0(16'b0011000100110011),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3571|_al_u3569  (
    .a({_al_u3569_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv }),
    .b({_al_u3570_o,_al_u3568_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({_al_u604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3571_o,_al_u3569_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*B))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~A*~(D*C*B))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0001010101010101),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3573|_al_u4282  (
    .a({_al_u3571_o,_al_u4281_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfjiu6 ,_al_u1296_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .f({_al_u3573_o,_al_u4282_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3575|_al_u3163  (
    .b({_al_u1344_o,open_n25902}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u1296_o,_al_u1344_o}),
    .f({_al_u3575_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3576|_al_u3220  (
    .b({_al_u1781_o,open_n25925}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u3575_o,_al_u677_o}),
    .f({_al_u3576_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C*~(~D*~A)))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C*~(~D*~A)))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000110001001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000110001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3577|_al_u1329  (
    .a({_al_u3574_o,open_n25950}),
    .b({_al_u3576_o,open_n25951}),
    .c({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u1329_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faoiu6 ,_al_u1329_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3578|_al_u3122  (
    .b({_al_u3122_o,open_n25978}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({_al_u1781_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u3578_o,_al_u3122_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*~A)))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~C*~(D*~(~B*~A)))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000100001111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000100001111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u357|_al_u6295  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12],_al_u6280_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13],_al_u6288_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14],_al_u5000_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15],_al_u6294_o}),
    .f({_al_u357_o,_al_u6295_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*A*~(D*~B))"),
    //.LUTF1("(~C*~B*~(D*A))"),
    //.LUTG0("(C*A*~(D*~B))"),
    //.LUTG1("(~C*~B*~(D*A))"),
    .INIT_LUTF0(16'b1000000010100000),
    .INIT_LUTF1(16'b0000000100000011),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b0000000100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3580|_al_u3579  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv }),
    .b({_al_u3578_o,_al_u2403_o}),
    .c({_al_u3579_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3580_o,_al_u3579_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3582|_al_u1635  (
    .b({_al_u678_o,open_n26049}),
    .c({_al_u679_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u1635_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u3582_o,_al_u1635_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3583|_al_u3128  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u3118_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u3583_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~D*~(~C*~B*~A))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000000011111110),
    .MODE("LOGIC"))
    \_al_u3585|_al_u3584  (
    .a({_al_u3582_o,_al_u678_o}),
    .b({_al_u3583_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u3584_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3585_o,_al_u3584_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+~(B)*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0101000000010101),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3586|_al_u3587  (
    .a({open_n26122,_al_u3586_o}),
    .b({open_n26123,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u3586_o,_al_u3587_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUT1("(~A*~(C*~(~D*B)))"),
    .INIT_LUT0(16'b0000010100001100),
    .INIT_LUT1(16'b0000010101000101),
    .MODE("LOGIC"))
    \_al_u3589|_al_u3588  (
    .a({_al_u3585_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .b({_al_u3587_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u2868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u3588_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0oiu6 ,_al_u3588_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u358|_al_u4859  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0],_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [0]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0]}),
    .f({_al_u358_o,_al_u4859_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~(C*B)*~(~D*A))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0011111100010101),
    .MODE("LOGIC"))
    \_al_u3590|_al_u1659  (
    .a({_al_u1659_o,open_n26188}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ifoiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({_al_u932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,_al_u1658_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdoiu6 ,_al_u1659_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(~D*~(A*~(C*B)))"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(~D*~(A*~(C*B)))"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b0000000011010101),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b0000000011010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3592|_al_u3591  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdoiu6 ,open_n26209}),
    .b({_al_u3591_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({_al_u1582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u3592_o,_al_u3591_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*A*~(D*~B))"),
    //.LUTF1("(~D*~(~C*B*A))"),
    //.LUTG0("(C*A*~(D*~B))"),
    //.LUTG1("(~D*~(~C*B*A))"),
    .INIT_LUTF0(16'b1000000010100000),
    .INIT_LUTF1(16'b0000000011110111),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b0000000011110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3593|_al_u3581  (
    .a({_al_u3581_o,_al_u3573_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0oiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Faoiu6 }),
    .c({_al_u3592_o,_al_u3580_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u3593_o,_al_u3581_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3595|_al_u1870  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aq2pw6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(B*A*~(D*~C))"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b1000000010001000),
    .MODE("LOGIC"))
    \_al_u3597|_al_u3596  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 }),
    .b({_al_u3596_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 }),
    .c({_al_u3120_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vmipw6 }),
    .f({_al_u3597_o,_al_u3596_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3598|_al_u3594  (
    .c({_al_u3593_o,_al_u1806_o}),
    .d({_al_u3132_o,_al_u3593_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 }));
  // ../RTL/cortexm0ds_logic.v(18745)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3599|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqlax6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u3597_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv }),
    .mi({open_n26340,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 }),
    .q({open_n26345,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] }));  // ../RTL/cortexm0ds_logic.v(18745)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u359|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6],open_n26346}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7],open_n26347}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n201 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u359_o,open_n26360}),
    .q({open_n26364,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(B*A*~(D*~C))"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b1000000010001000),
    .MODE("LOGIC"))
    \_al_u3601|_al_u3600  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpniu6 }),
    .c({_al_u3120_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 }),
    .f({_al_u3601_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Inniu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(B*A*~(D*~C))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(B*A*~(D*~C))"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000000010001000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3603|_al_u3121  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Crniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqniu6 ,_al_u3120_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yoniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 }),
    .f({_al_u3603_o,_al_u3121_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u360|_al_u4625  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2],_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [3]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3]}),
    .f({_al_u360_o,_al_u4625_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*C*B))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b1010101000101010),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u3610|_al_u3609  (
    .a({open_n26429,_al_u3608_o}),
    .b({_al_u3609_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({_al_u2365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3610_o,_al_u3609_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(C*~(~B*~(~D*A)))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1100000011100000),
    .MODE("LOGIC"))
    \_al_u3612|_al_u3611  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv }),
    .b({_al_u3611_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 }),
    .c({_al_u1582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3612_o,_al_u3611_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*C*A))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(~B*~(D*C*A))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0001001100110011),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0001001100110011),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3615|_al_u3614  (
    .a({_al_u3157_o,_al_u3110_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({_al_u3614_o,_al_u2829_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3615_o,_al_u3614_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(A*(B@(~D*C)))"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(A*(B@(~D*C)))"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1000100000101000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b1000100000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3616|_al_u3652  (
    .a({_al_u3215_o,_al_u3215_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro1ju6 ,_al_u3652_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(~C*A))"),
    //.LUT1("(C*B*~(D*A))"),
    .INIT_LUT0(16'b0000000000110001),
    .INIT_LUT1(16'b0100000011000000),
    .MODE("LOGIC"))
    \_al_u3617|_al_u6252  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 }),
    .b({_al_u3613_o,_al_u6251_o}),
    .c({_al_u3615_o,_al_u2380_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro1ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({_al_u3617_o,_al_u6252_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000011101010),
    .MODE("LOGIC"))
    \_al_u3619|_al_u3618  (
    .a({_al_u3618_o,open_n26538}),
    .b({_al_u681_o,_al_u607_o}),
    .c({_al_u2829_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jr1ju6_lutinv ,_al_u3618_o}));
  // ../RTL/cortexm0ds_logic.v(17470)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(~B*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~(~D*C)*~(~B*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110100001101),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1101110100001101),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3620|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6_reg  (
    .a({_al_u3610_o,_al_u3620_o}),
    .b({_al_u3617_o,_al_u3622_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jr1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1342_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 }),
    .f({_al_u3620_o,open_n26577}),
    .q({open_n26581,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 }));  // ../RTL/cortexm0ds_logic.v(17470)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3622|_al_u3621  (
    .b({_al_u3110_o,_al_u3109_o}),
    .c({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u3621_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv }),
    .f({_al_u3622_o,_al_u3621_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u3625|_al_u930  (
    .a({_al_u2364_o,open_n26608}),
    .b({_al_u930_o,open_n26609}),
    .c({_al_u2764_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u3625_o,_al_u930_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(B*~A*~(~D*C))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0100010000000100),
    .MODE("LOGIC"))
    \_al_u3626|_al_u3624  (
    .a({_al_u3624_o,open_n26630}),
    .b({_al_u3625_o,open_n26631}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,_al_u909_o}),
    .f({_al_u3626_o,_al_u3624_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u3630|_al_u3629  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 ,open_n26652}),
    .b({_al_u3629_o,open_n26653}),
    .c({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .f({_al_u3630_o,_al_u3629_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(D*C))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(~B*~A*~(D*C))"),
    //.LUTG1("(D*C*~B*A)"),
    .INIT_LUTF0(16'b0000000100010001),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0000000100010001),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3631|_al_u3628  (
    .a({_al_u3627_o,_al_u2758_o}),
    .b({_al_u3189_o,_al_u1583_o}),
    .c({_al_u3628_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .d({_al_u3630_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3631_o,_al_u3628_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3633|_al_u3632  (
    .b({_al_u3632_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bziiu6_lutinv ,_al_u606_o}),
    .f({_al_u3633_o,_al_u3632_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*A*~(D*B))"),
    //.LUT1("(B*A*~(D*~C))"),
    .INIT_LUT0(16'b0000001000001010),
    .INIT_LUT1(16'b1000000010001000),
    .MODE("LOGIC"))
    \_al_u3636|_al_u3635  (
    .a({_al_u3631_o,_al_u3633_o}),
    .b({_al_u3635_o,_al_u1812_o}),
    .c({_al_u1643_o,_al_u3634_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3636_o,_al_u3635_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~D*~C*B))"),
    //.LUT1("(~D*~C*B*A)"),
    .INIT_LUT0(16'b0101010101010001),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"))
    \_al_u3637|_al_u3638  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 ,_al_u3637_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3637_o,_al_u3638_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*~A)"),
    //.LUT1("(B*~A*~(~D*~C))"),
    .INIT_LUT0(16'b0000010000000000),
    .INIT_LUT1(16'b0100010001000000),
    .MODE("LOGIC"))
    \_al_u3640|_al_u3639  (
    .a({_al_u3638_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .b({_al_u3639_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .f({_al_u3640_o,_al_u3639_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~C)*~(~B*A))"),
    //.LUTF1("(~C*~A*~(D*~B))"),
    //.LUTG0("(~(D*~C)*~(~B*A))"),
    //.LUTG1("(~C*~A*~(D*~B))"),
    .INIT_LUTF0(16'b1101000011011101),
    .INIT_LUTF1(16'b0000010000000101),
    .INIT_LUTG0(16'b1101000011011101),
    .INIT_LUTG1(16'b0000010000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3642|_al_u3641  (
    .a({_al_u1802_o,_al_u1342_o}),
    .b({_al_u3641_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ,_al_u3641_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~C*B))"),
    //.LUTF1("(C*A*~(D*~B))"),
    //.LUTG0("(A*~(~D*~C*B))"),
    //.LUTG1("(C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1010101010100010),
    .INIT_LUTF1(16'b1000000010100000),
    .INIT_LUTG0(16'b1010101010100010),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3643|_al_u3646  (
    .a({_al_u3636_o,_al_u3643_o}),
    .b({_al_u3640_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u3643_o,_al_u3646_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(A*~(D*~C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b1010001010101010),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1010001010101010),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3647|_al_u3648  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ,_al_u3647_o}),
    .b({_al_u2364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3647_o,_al_u3648_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u3649|_al_u3215  (
    .b({_al_u912_o,open_n26858}),
    .c({_al_u3215_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({_al_u3648_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u3649_o,_al_u3215_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(~B*~(D*~(~C*~A)))"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b0000000100110011),
    .MODE("LOGIC"))
    \_al_u3651|_al_u3650  (
    .a({_al_u2380_o,open_n26879}),
    .b({_al_u3650_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ,_al_u3650_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(A*~(C)*~(D)+~(A)*C*D))"),
    //.LUT1("(C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000000001000),
    .INIT_LUT1(16'b1111000011010000),
    .MODE("LOGIC"))
    \_al_u3654|_al_u3653  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .b({_al_u3652_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({_al_u2364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({_al_u3653_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3654_o,_al_u3653_o}));
  // ../RTL/cortexm0ds_logic.v(17277)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(A*~(D*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111011100000101),
    .INIT_LUT1(16'b0000100010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3655|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6_reg  (
    .a({_al_u3646_o,_al_u3655_o}),
    .b({_al_u3649_o,_al_u3659_o}),
    .c({_al_u3654_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3655_o,open_n26933}),
    .q({open_n26937,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }));  // ../RTL/cortexm0ds_logic.v(17277)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~B*~(C*A)))"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .INIT_LUT0(16'b0000000011101100),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"))
    \_al_u3659|_al_u3658  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv ,_al_u607_o}),
    .b({_al_u3657_o,_al_u2813_o}),
    .c({_al_u3658_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u3094_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3659_o,_al_u3658_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*~C*B))"),
    //.LUT1("(~A*~(D*~C*B))"),
    .INIT_LUT0(16'b0101000101010101),
    .INIT_LUT1(16'b0101000101010101),
    .MODE("LOGIC"))
    \_al_u3663|_al_u3662  (
    .a({_al_u3661_o,_al_u2365_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({_al_u3662_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3663_o,_al_u3662_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3664|_al_u3232  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujjiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 }),
    .f({_al_u3664_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~B*A*~(~D*C))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~B*A*~(~D*C))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0010001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3665|_al_u3645  (
    .a({_al_u3663_o,open_n27004}),
    .b({_al_u3664_o,open_n27005}),
    .c({_al_u2847_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv }),
    .f({_al_u3665_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3666|_al_u2825  (
    .b({open_n27032,_al_u2824_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yecpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({_al_u3629_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 }),
    .f({_al_u3666_o,_al_u2825_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3667|_al_u3236  (
    .b({open_n27059,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u3236_o,_al_u609_o}),
    .f({_al_u3667_o,_al_u3236_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(~D*A))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0011111100010101),
    .MODE("LOGIC"))
    \_al_u3669|_al_u2844  (
    .a({_al_u3187_o,open_n27080}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv ,open_n27081}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3669_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K49ow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*A*~(~D*C))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0010001000000010),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u3672|_al_u3670  (
    .a({open_n27102,_al_u909_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({_al_u1662_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u3670_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3672_o,_al_u3670_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3673|_al_u3668  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T41ju6 ,_al_u3666_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U99ow6 ,_al_u3667_o}),
    .c({_al_u3669_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({_al_u3672_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u3673_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U99ow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~B*A)"),
    //.LUT1("(A*~(~C*~(D*B)))"),
    .INIT_LUT0(16'b0000000000100000),
    .INIT_LUT1(16'b1010100010100000),
    .MODE("LOGIC"))
    \_al_u3675|_al_u3674  (
    .a({_al_u3109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u3674_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3675_o,_al_u3674_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(A*~(C*~B)))"),
    //.LUTF1("(A*~(~B*~(~D*C)))"),
    //.LUTG0("(D*~(A*~(C*~B)))"),
    //.LUTG1("(A*~(~B*~(~D*C)))"),
    .INIT_LUTF0(16'b0111010100000000),
    .INIT_LUTF1(16'b1000100010101000),
    .INIT_LUTG0(16'b0111010100000000),
    .INIT_LUTG1(16'b1000100010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3677|_al_u3676  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .b({_al_u2772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kb9ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3677_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kb9ow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*~A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~D*C*B*~A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b0000000001000000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000001000000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3678|_al_u3834  (
    .a({_al_u3665_o,_al_u3827_o}),
    .b({_al_u3673_o,_al_u3830_o}),
    .c({_al_u3675_o,_al_u3832_o}),
    .d({_al_u3677_o,_al_u3833_o}),
    .f({_al_u3678_o,_al_u3834_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~A*~(D*B))"),
    //.LUTF1("(B*A*~(~D*~C))"),
    //.LUTG0("(~C*~A*~(D*B))"),
    //.LUTG1("(B*A*~(~D*~C))"),
    .INIT_LUTF0(16'b0000000100000101),
    .INIT_LUTF1(16'b1000100010000000),
    .INIT_LUTG0(16'b0000000100000101),
    .INIT_LUTG1(16'b1000100010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3679|_al_u3234  (
    .a({_al_u3214_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3679_o,_al_u3234_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3680|_al_u2369  (
    .c({_al_u2369_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u3680_o,_al_u2369_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    //.LUT1("(B*~(A*~(~D*C)))"),
    .INIT_LUT0(16'b0010001000000011),
    .INIT_LUT1(16'b0100010011000100),
    .MODE("LOGIC"))
    \_al_u3684|_al_u3683  (
    .a({_al_u3681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .b({_al_u2770_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u3683_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3684_o,_al_u3683_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*B*C*D)"),
    //.LUT1("(A*~(~B*~(~D*C)))"),
    .INIT_LUT0(16'b1000110111111011),
    .INIT_LUT1(16'b1000100010101000),
    .MODE("LOGIC"))
    \_al_u3686|_al_u3685  (
    .a({_al_u2386_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .b({_al_u2764_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh9ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3686_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh9ow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3689|_al_u2371  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({_al_u2371_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ,_al_u2371_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"))
    \_al_u3691|_al_u3690  (
    .a({_al_u912_o,open_n27331}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ,open_n27332}),
    .c({_al_u3690_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u696_o,_al_u1344_o}),
    .f({_al_u3691_o,_al_u3690_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A*~(~C*B)))"),
    //.LUT1("(D*~C*~B*~A)"),
    .INIT_LUT0(16'b0101110100000000),
    .INIT_LUT1(16'b0000000100000000),
    .MODE("LOGIC"))
    \_al_u3692|_al_u3688  (
    .a({_al_u3684_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Io9ow6 }),
    .b({_al_u3686_o,_al_u1367_o}),
    .c({_al_u3688_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u3691_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3692_o,_al_u3688_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    //.LUTF1("(C*~(~B*~(D*~A)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    //.LUTG1("(C*~(~B*~(D*~A)))"),
    .INIT_LUTF0(16'b0000110011110101),
    .INIT_LUTF1(16'b1101000011000000),
    .INIT_LUTG0(16'b0000110011110101),
    .INIT_LUTG1(16'b1101000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3694|_al_u3693  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ,_al_u1643_o}),
    .b({_al_u3693_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({_al_u1806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u3694_o,_al_u3693_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*A*~(~D*~B))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000101000001000),
    .MODE("LOGIC"))
    \_al_u3695|_al_u3095  (
    .a({_al_u3678_o,open_n27397}),
    .b({_al_u3692_o,open_n27398}),
    .c({_al_u3694_o,_al_u3094_o}),
    .d({_al_u1812_o,_al_u1812_o}),
    .f({_al_u3695_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17741)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(~B*A))"),
    //.LUTF1("(D*~A*~(~C*~B))"),
    //.LUTG0("(~(~D*C)*~(~B*A))"),
    //.LUTG1("(D*~A*~(~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110100001101),
    .INIT_LUTF1(16'b0101010000000000),
    .INIT_LUTG0(16'b1101110100001101),
    .INIT_LUTG1(16'b0101010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3697|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6_reg  (
    .a({_al_u3696_o,_al_u3695_o}),
    .b({_al_u607_o,_al_u3697_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3697_o,open_n27436}),
    .q({open_n27440,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }));  // ../RTL/cortexm0ds_logic.v(17741)
  // ../RTL/cortexm0ds_logic.v(19131)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3699|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ,open_n27441}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ,open_n27442}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ,_al_u2506_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({open_n27453,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3699_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n127 }),
    .q({open_n27457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 }));  // ../RTL/cortexm0ds_logic.v(19131)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3700|_al_u3987  (
    .a({_al_u3271_o,open_n27458}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 }),
    .f({_al_u3700_o,_al_u3987_o}));
  // ../RTL/cortexm0ds_logic.v(19707)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3701|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ,open_n27483}),
    .b({_al_u3446_o,\u_cmsdk_mcu/sram_hrdata [30]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ,\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ,\u_cmsdk_mcu/HWDATA [30]}),
    .mi({open_n27487,\u_cmsdk_mcu/HWDATA [30]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3701_o,\u_cmsdk_mcu/u_ahb_ram/n13 [30]}),
    .q({open_n27502,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 }));  // ../RTL/cortexm0ds_logic.v(19707)
  // ../RTL/cortexm0ds_logic.v(19077)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3702|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6_reg  (
    .a({_al_u3454_o,open_n27503}),
    .b({_al_u3463_o,open_n27504}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ,_al_u2518_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({open_n27515,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3702_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n127 }),
    .q({open_n27519,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 }));  // ../RTL/cortexm0ds_logic.v(19077)
  // ../RTL/cortexm0ds_logic.v(19587)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3704|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ,open_n27520}),
    .b({_al_u3520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ,\u_cmsdk_mcu/HWDATA [30]}),
    .mi({open_n27524,\u_cmsdk_mcu/HWDATA [30]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3704_o,_al_u3517_o}),
    .q({open_n27539,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 }));  // ../RTL/cortexm0ds_logic.v(19587)
  // ../RTL/cortexm0ds_logic.v(19653)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*D))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("~(~C*~(B*D))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011110000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1111110011110000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3705|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6_reg  (
    .a({_al_u3703_o,open_n27540}),
    .b({_al_u3704_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write1 }),
    .c({_al_u3530_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [14]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({open_n27544,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3705_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n299 }),
    .q({open_n27559,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 }));  // ../RTL/cortexm0ds_logic.v(19653)
  // ../RTL/cortexm0ds_logic.v(20118)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3706|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv ,open_n27560}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odfiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ,_al_u3274_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3706_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4phu6 }),
    .q({open_n27581,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 }));  // ../RTL/cortexm0ds_logic.v(20118)
  // ../RTL/cortexm0ds_logic.v(19005)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3707|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6_reg  (
    .a({_al_u3281_o,open_n27582}),
    .b({_al_u3479_o,open_n27583}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ,_al_u2514_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({open_n27587,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3707_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n217 }),
    .q({open_n27602,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 }));  // ../RTL/cortexm0ds_logic.v(19005)
  // ../RTL/cortexm0ds_logic.v(19341)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3708|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6_reg  (
    .a({_al_u3372_o,open_n27603}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ,_al_u3352_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3708_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2phu6 }),
    .q({open_n27624,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 }));  // ../RTL/cortexm0ds_logic.v(19341)
  // ../RTL/cortexm0ds_logic.v(19605)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3709|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ,open_n27625}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ,open_n27626}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ,_al_u2516_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({open_n27637,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3709_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n172 }),
    .q({open_n27641,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 }));  // ../RTL/cortexm0ds_logic.v(19605)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~((~C*~B))*~(D)+A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000001111111110),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u370|_al_u364  (
    .a({open_n27642,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]}),
    .b({open_n27643,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3:2]),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]}),
    .f({_al_u370_o,_al_u364_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3710|_al_u3722  (
    .a({_al_u3706_o,_al_u3705_o}),
    .b({_al_u3707_o,_al_u3710_o}),
    .c({_al_u3708_o,_al_u3716_o}),
    .d({_al_u3709_o,_al_u3721_o}),
    .f({_al_u3710_o,_al_u3722_o}));
  // ../RTL/cortexm0ds_logic.v(19317)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3711|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ,open_n27688}),
    .b({_al_u3443_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ,_al_u3345_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isbpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2phu6 }),
    .q({open_n27705,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 }));  // ../RTL/cortexm0ds_logic.v(19317)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"))
    \_al_u3712|_al_u3349  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ,open_n27708}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8row6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljbpw6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3714|_al_u3946  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ,open_n27729}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2cpw6 ,_al_u3946_o}));
  // ../RTL/cortexm0ds_logic.v(19689)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3715|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6_reg  (
    .a({_al_u3468_o,open_n27754}),
    .b({_al_u3350_o,open_n27755}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ,_al_u2520_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({open_n27759,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3715_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n82 }),
    .q({open_n27774,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 }));  // ../RTL/cortexm0ds_logic.v(19689)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3716|_al_u3713  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isbpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 }),
    .b({_al_u3713_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2cpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 }),
    .d({_al_u3715_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 }),
    .f({_al_u3716_o,_al_u3713_o}));
  // ../RTL/cortexm0ds_logic.v(17206)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~A*~(D*~C))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~A*~(D*~C))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111110111011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1011111110111011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3717|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 ,_al_u2121_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ,_al_u2128_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 ,_al_u2272_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3717_o,\u_cmsdk_mcu/HWDATA [30]}),
    .q({open_n27818,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 }));  // ../RTL/cortexm0ds_logic.v(17206)
  // ../RTL/cortexm0ds_logic.v(19920)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3718|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6_reg  (
    .a({_al_u3335_o,open_n27819}),
    .b({_al_u3343_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ,_al_u3343_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ,_al_u3342_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3718_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V4phu6 }),
    .q({open_n27840,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 }));  // ../RTL/cortexm0ds_logic.v(19920)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u3720|_al_u3981  (
    .a({_al_u3489_o,open_n27841}),
    .b({_al_u3515_o,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 ,_al_u3489_o}),
    .f({_al_u3720_o,_al_u3981_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u3721|_al_u3719  (
    .a({_al_u3717_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv }),
    .b({_al_u3718_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv }),
    .c({_al_u3719_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 }),
    .d({_al_u3720_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 }),
    .f({_al_u3721_o,_al_u3719_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3723|_al_u6585  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 }),
    .d({_al_u3722_o,_al_u6333_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vwapw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffrow6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(19329)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3724|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6_reg  (
    .a({_al_u3343_o,open_n27910}),
    .b({_al_u3350_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ,_al_u3350_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ,_al_u3348_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3724_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K2phu6 }),
    .q({open_n27927,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 }));  // ../RTL/cortexm0ds_logic.v(19329)
  // ../RTL/cortexm0ds_logic.v(19713)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3725|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv ,open_n27928}),
    .b({_al_u3446_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ,\u_cmsdk_mcu/HWDATA [31]}),
    .mi({open_n27939,\u_cmsdk_mcu/HWDATA [31]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3725_o,_al_u3522_o}),
    .q({open_n27943,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 }));  // ../RTL/cortexm0ds_logic.v(19713)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3726|_al_u3966  (
    .a({_al_u3463_o,open_n27944}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ,_al_u3463_o}),
    .f({_al_u3726_o,_al_u3966_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u3727|_al_u3926  (
    .a({_al_u3443_o,open_n27969}),
    .b({_al_u3520_o,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ,_al_u3520_o}),
    .f({_al_u3727_o,_al_u3926_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3728|_al_u6432  (
    .a({_al_u3724_o,open_n27990}),
    .b({_al_u3725_o,open_n27991}),
    .c({_al_u3726_o,_al_u6423_o}),
    .d({_al_u3727_o,_al_u6421_o}),
    .f({_al_u3728_o,_al_u6432_o}));
  // ../RTL/cortexm0ds_logic.v(19677)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*~A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*~A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010101000111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0010101000111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3729|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ,_al_u3874_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ,\u_cmsdk_mcu/HWDATA [31]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 }),
    .mi({open_n28019,\u_cmsdk_mcu/HWDATA [31]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3729_o,_al_u3875_o}),
    .q({open_n28034,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 }));  // ../RTL/cortexm0ds_logic.v(19677)
  // ../RTL/cortexm0ds_logic.v(20266)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~A*~(D*C*~B))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~A*~(D*C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0100010101010101),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0100010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u372|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6_reg  (
    .a({XTAL1_wire,open_n28035}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usaiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3row6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 ,_al_u6596_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({XTAL2_pad,open_n28052}),
    .q({open_n28056,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cokbx6 }));  // ../RTL/cortexm0ds_logic.v(20266)
  // ../RTL/cortexm0ds_logic.v(19659)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3730|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6_reg  (
    .a({_al_u3728_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 }),
    .b({_al_u3729_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 }),
    .c({_al_u3530_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 }),
    .mi({open_n28060,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3730_o,_al_u6690_o}),
    .q({open_n28075,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 }));  // ../RTL/cortexm0ds_logic.v(19659)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u3731|_al_u5386  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 }),
    .f({_al_u3731_o,_al_u5386_o}));
  // ../RTL/cortexm0ds_logic.v(19629)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3732|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dagiu6_lutinv ,open_n28096}),
    .b({_al_u3468_o,\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ,\u_cmsdk_mcu/flash_hrdata [31]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ,\u_cmsdk_mcu/HWDATA [31]}),
    .mi({open_n28107,\u_cmsdk_mcu/HWDATA [31]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3732_o,\u_cmsdk_mcu/u_ahb_rom/n13 [31]}),
    .q({open_n28111,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 }));  // ../RTL/cortexm0ds_logic.v(19629)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3735|_al_u3733  (
    .a({_al_u3731_o,_al_u3271_o}),
    .b({_al_u3732_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 }),
    .c({_al_u3733_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 }),
    .d({_al_u3734_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 }),
    .f({_al_u3735_o,_al_u3733_o}));
  // ../RTL/cortexm0ds_logic.v(20200)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3737|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv ,open_n28136}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eegiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ,_al_u3286_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3bpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwdpw6 }),
    .q({open_n28153,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 }));  // ../RTL/cortexm0ds_logic.v(20200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3738|_al_u5382  (
    .a({_al_u3489_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ,_al_u546_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 }),
    .f({_al_u3738_o,_al_u5382_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u3739|_al_u3975  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 ,open_n28178}),
    .b({_al_u3479_o,_al_u3925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ,_al_u3479_o}),
    .f({_al_u3739_o,_al_u3975_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3740|_al_u3736  (
    .a({_al_u3736_o,_al_u3335_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3bpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ajgiu6 }),
    .c({_al_u3738_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 }),
    .d({_al_u3739_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 }),
    .f({_al_u3740_o,_al_u3736_o}));
  // ../RTL/cortexm0ds_logic.v(19053)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3741|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6_reg  (
    .a({_al_u3372_o,open_n28223}),
    .b({_al_u3454_o,\u_cmsdk_mcu/HWDATA [31]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 ,_al_u2725_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ,_al_u3780_o}),
    .mi({open_n28227,\u_cmsdk_mcu/HWDATA [31]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3741_o,_al_u3781_o}),
    .q({open_n28242,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 }));  // ../RTL/cortexm0ds_logic.v(19053)
  // ../RTL/cortexm0ds_logic.v(19701)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3742|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ,open_n28243}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3giu6 ,\u_cmsdk_mcu/sram_hrdata [23]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ,\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ,\u_cmsdk_mcu/HWDATA [23]}),
    .mi({open_n28247,\u_cmsdk_mcu/HWDATA [23]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3742_o,\u_cmsdk_mcu/u_ahb_ram/n13 [23]}),
    .q({open_n28262,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 }));  // ../RTL/cortexm0ds_logic.v(19701)
  // ../RTL/cortexm0ds_logic.v(19035)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3743|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6_reg  (
    .a({_al_u3281_o,open_n28263}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ,open_n28264}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ,\u_cmsdk_mcu/HWDATA [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3743_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 }),
    .q({open_n28284,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 }));  // ../RTL/cortexm0ds_logic.v(19035)
  // ../RTL/cortexm0ds_logic.v(19563)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3744|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ,open_n28285}),
    .b({_al_u3515_o,open_n28286}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ,_al_u2476_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n28297,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3744_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n248 }),
    .q({open_n28301,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 }));  // ../RTL/cortexm0ds_logic.v(19563)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3745|_al_u6492  (
    .a({_al_u3741_o,open_n28302}),
    .b({_al_u3742_o,open_n28303}),
    .c({_al_u3743_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 }),
    .d({_al_u3744_o,_al_u6464_o}),
    .f({_al_u3745_o,_al_u6492_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u3746|_al_u6336  (
    .a({_al_u3730_o,open_n28328}),
    .b({_al_u3735_o,open_n28329}),
    .c({_al_u3740_o,_al_u6335_o}),
    .d({_al_u3745_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ,_al_u6336_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3748|_al_u3380  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejbpw6 }),
    .f({_al_u3748_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhgiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3749|_al_u3747  (
    .b({_al_u3748_o,open_n28376}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uybpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmbpw6 }),
    .d({_al_u3747_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 }),
    .f({_al_u3749_o,_al_u3747_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(~C*(~(A)*B*~(D)+~(A)*~(B)*D+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0000110100000100),
    .MODE("LOGIC"))
    \_al_u3750|_al_u3751  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vwapw6 ,open_n28401}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 }),
    .c({_al_u3749_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ,_al_u3750_o}),
    .f({_al_u3750_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3752|_al_u3753  (
    .b({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utgiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utgiu6 ,_al_u3753_o}));
  // ../RTL/cortexm0ds_logic.v(19695)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(A*~(~B*~(D*C)))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(A*~(~B*~(D*C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1010100010001000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1010100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3755|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ,open_n28444}),
    .b({_al_u3753_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 }),
    .c({_al_u3754_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u3124_o,_al_u3755_o}),
    .mi({open_n28448,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3755_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 }),
    .q({open_n28463,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 }));  // ../RTL/cortexm0ds_logic.v(19695)
  // ../RTL/cortexm0ds_logic.v(18959)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3756|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 }),
    .mi({open_n28467,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ,_al_u6692_o}),
    .q({open_n28483,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9xax6 }));  // ../RTL/cortexm0ds_logic.v(18959)
  // ../RTL/cortexm0ds_logic.v(18079)
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(D*~(C*B)))"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("~(A*~(D*~(C*B)))"),
    //.LUTG1("(C*~(B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111101010101),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b0111111101010101),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3758|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6_reg  (
    .a({open_n28484,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrgiu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrgiu6 ,_al_u3758_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3758_o,open_n28502}),
    .q({open_n28506,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 }));  // ../RTL/cortexm0ds_logic.v(18079)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u375|_al_u503  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .d({_al_u374_o,_al_u374_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3760|_al_u3767  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv }),
    .d({_al_u3597_o,_al_u3597_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3762|_al_u3764  (
    .c({_al_u3603_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkniu6_lutinv }),
    .d({_al_u3601_o,_al_u3597_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17851)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3769|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hoxpw6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 }),
    .mi({open_n28603,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({_al_u3769_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 }),
    .q({open_n28608,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[10] }));  // ../RTL/cortexm0ds_logic.v(17851)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*~C*~B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000001000000000),
    .MODE("LOGIC"))
    \_al_u376|_al_u5022  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vowiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }));
  // ../RTL/cortexm0ds_logic.v(18893)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3771|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewtax6_reg  (
    .c({_al_u3603_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u3601_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhniu6_lutinv }),
    .mi({open_n28643,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 }),
    .q({open_n28648,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[10] }));  // ../RTL/cortexm0ds_logic.v(18893)
  // ../RTL/cortexm0ds_logic.v(20272)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D*~(C*~A)))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(D*~(C*~A)))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1011111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3777|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqkbx6_reg  (
    .a({open_n28649,_al_u3776_o}),
    .b({_al_u1676_o,_al_u3777_o}),
    .c({\u_cmsdk_mcu/dbg_swdo_en ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1253_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u3777_o,open_n28667}),
    .q({open_n28671,\u_cmsdk_mcu/dbg_swdo_en }));  // ../RTL/cortexm0ds_logic.v(20272)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3779|_al_u3137  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .f({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000110011111100),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3782|_al_u2735  (
    .b({_al_u2733_o,\u_cmsdk_mcu/sram_hrdata [28]}),
    .c({_al_u2741_o,\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}),
    .d({_al_u2729_o,_al_u2733_o}),
    .f({_al_u3782_o,\u_cmsdk_mcu/u_ahb_ram/n13 [28]}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3785|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b18  (
    .a({_al_u3781_o,\u_cmsdk_mcu/HWDATA [18]}),
    .b({_al_u3782_o,\u_cmsdk_mcu/HWDATA [19]}),
    .c({_al_u3783_o,\u_cmsdk_mcu/HWDATA [20]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({_al_u3784_o,\u_cmsdk_mcu/HWDATA [21]}),
    .mi({open_n28728,\u_cmsdk_mcu/HWDATA [18]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 ,_al_u3784_o}),
    .q({open_n28732,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [18]}));  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*B))"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~A*~(D*C*B))"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b0001010101010101),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3788|_al_u3787  (
    .a({open_n28733,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G1aow6 }),
    .b({_al_u3787_o,_al_u607_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u3788_o,_al_u3787_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~B*~(~D*A)))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~C*~(~B*~(~D*A)))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000110000001110),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000110000001110),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3789|_al_u3157  (
    .a({open_n28758,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .b({_al_u3156_o,_al_u3156_o}),
    .c({_al_u2392_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u3789_o,_al_u3157_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u3790|_al_u3797  (
    .a({open_n28783,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 }),
    .b({_al_u1297_o,_al_u3788_o}),
    .c({_al_u606_o,_al_u3790_o}),
    .d({_al_u3789_o,_al_u3796_o}),
    .f({_al_u3790_o,_al_u3797_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3791|_al_u697  (
    .a({_al_u697_o,_al_u695_o}),
    .b({_al_u3159_o,_al_u696_o}),
    .c({_al_u609_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3791_o,_al_u697_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u3794|_al_u3793  (
    .a({open_n28828,_al_u696_o}),
    .b({_al_u3793_o,_al_u2392_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv }),
    .d({_al_u3624_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3794_o,_al_u3793_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*~A)"),
    //.LUT1("(~D*C*~B*A)"),
    .INIT_LUT0(16'b0000000001000000),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u3796|_al_u3795  (
    .a({_al_u3791_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .b({_al_u3792_o,_al_u1266_o}),
    .c({_al_u3794_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u3795_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u3796_o,_al_u3795_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(D*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1010100011111100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u379|_al_u557  (
    .a({open_n28869,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n31 }),
    .b({open_n28870,uart0_txen_pad}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [0]}),
    .f({_al_u379_o,_al_u557_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~B*~(D*C)))"),
    //.LUT1("(D*~C*~B*~A)"),
    .INIT_LUT0(16'b1010100010001000),
    .INIT_LUT1(16'b0000000100000000),
    .MODE("LOGIC"))
    \_al_u3801|_al_u3800  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u3800_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u3801_o,_al_u3800_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~((D*B))*~(C)+A*(D*B)*~(C)+~(A)*(D*B)*C+A*(D*B)*C)"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("~(A*~((D*B))*~(C)+A*(D*B)*~(C)+~(A)*(D*B)*C+A*(D*B)*C)"),
    //.LUTG1("(~A*~(D*C*B))"),
    .INIT_LUTF0(16'b0011010111110101),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b0011010111110101),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3802|_al_u3798  (
    .a({_al_u3797_o,_al_u682_o}),
    .b({_al_u3798_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .c({_al_u3799_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u3801_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u3798_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3803|_al_u2801  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .f({_al_u3803_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*~A*~(D*B))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000100000101),
    .MODE("LOGIC"))
    \_al_u3805|_al_u3804  (
    .a({_al_u3803_o,open_n28959}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ,_al_u2813_o}),
    .c({_al_u3804_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,_al_u604_o}),
    .f({_al_u3805_o,_al_u3804_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"))
    \_al_u3806|_al_u2410  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ,open_n28980}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ,open_n28981}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u3806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~A*~(~D*C*B))"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~A*~(~D*C*B))"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0101010100010101),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0101010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3808|_al_u3807  (
    .a({_al_u3797_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .b({_al_u3805_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({_al_u3806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u3807_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u3808_o,_al_u3807_o}));
  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u380|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b2  (
    .a({_al_u379_o,open_n29026}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0],open_n29027}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ,open_n29040}),
    .q({open_n29044,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [2]}));  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3810|_al_u2753  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv }),
    .f({_al_u3810_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~(D*~A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*B*~(D*~A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000100000001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000100000001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3811|_al_u4044  (
    .a({open_n29073,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9aiu6 }),
    .b({open_n29074,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({_al_u3811_o,_al_u4044_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~(C*~B)*~(D*A))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~(C*~B)*~(D*A))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0100010111001111),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0100010111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3813|_al_u3812  (
    .a({_al_u3810_o,_al_u1812_o}),
    .b({_al_u3812_o,_al_u2380_o}),
    .c({_al_u903_o,_al_u3811_o}),
    .d({_al_u1342_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({_al_u3813_o,_al_u3812_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u3815|_al_u3814  (
    .a({open_n29123,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv }),
    .b({_al_u1782_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({_al_u3814_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3815_o,_al_u3814_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u3818|_al_u3817  (
    .a({_al_u3815_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .b({_al_u3816_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({_al_u3817_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3818_o,_al_u3817_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(~B*~(~D*~C*A))"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(~B*~(~D*~C*A))"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0011001100110001),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0011001100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3820|_al_u3150  (
    .a({_al_u3629_o,open_n29164}),
    .b({_al_u3819_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u3150_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 }),
    .f({_al_u3820_o,_al_u3150_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))"),
    //.LUTF1("(B*~(D*~C*A))"),
    //.LUTG0("(A*(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))"),
    //.LUTG1("(B*~(D*~C*A))"),
    .INIT_LUTF0(16'b1000100000001010),
    .INIT_LUTF1(16'b1100010011001100),
    .INIT_LUTG0(16'b1000100000001010),
    .INIT_LUTG1(16'b1100010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3821|_al_u3559  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 }),
    .b({_al_u3820_o,_al_u1266_o}),
    .c({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btoiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3821_o,_al_u3559_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(D*~A))"),
    //.LUT1("(A*~(D*C*B))"),
    .INIT_LUT0(16'b1000000011000000),
    .INIT_LUT1(16'b0010101010101010),
    .MODE("LOGIC"))
    \_al_u3823|_al_u3822  (
    .a({_al_u3822_o,_al_u3813_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv ,_al_u3818_o}),
    .c({_al_u2754_o,_al_u3821_o}),
    .d({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u3823_o,_al_u3822_o}));
  // ../RTL/cortexm0ds_logic.v(17518)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(~B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(~D*C)*~(~B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110100001101),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1101110100001101),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3825|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6_reg  (
    .a({open_n29233,_al_u3825_o}),
    .b({_al_u3824_o,_al_u3849_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u3823_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3825_o,open_n29251}),
    .q({open_n29255,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }));  // ../RTL/cortexm0ds_logic.v(17518)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3827|_al_u3826  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ,open_n29258}),
    .c({_al_u3826_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u1643_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u3827_o,_al_u3826_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~A*~(B*~(~D*~C)))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0001000100010101),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0001000100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3828|_al_u2775  (
    .a({_al_u2772_o,open_n29283}),
    .b({_al_u2364_o,open_n29284}),
    .c({_al_u2764_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc6ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*A*~(C*~B))"),
    //.LUT1("(~C*A*~(D*B))"),
    .INIT_LUT0(16'b0000000010001010),
    .INIT_LUT1(16'b0000001000001010),
    .MODE("LOGIC"))
    \_al_u3830|_al_u3829  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc6ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .b({_al_u1799_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 }),
    .c({_al_u3829_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u3830_o,_al_u3829_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~(D*B)*~(~C*A))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~(D*B)*~(~C*A))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0011000111110101),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0011000111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3832|_al_u3831  (
    .a({_al_u3754_o,open_n29329}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ,open_n29330}),
    .c({_al_u1813_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u3831_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u3832_o,_al_u3831_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3833|_al_u4379  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ,_al_u3246_o}),
    .f({_al_u3833_o,_al_u4379_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~A*~(D*B)))"),
    //.LUT1("(A*~(D*C*B))"),
    .INIT_LUT0(16'b0000111000001010),
    .INIT_LUT1(16'b0010101010101010),
    .MODE("LOGIC"))
    \_al_u3836|_al_u3835  (
    .a({_al_u3834_o,_al_u604_o}),
    .b({_al_u3109_o,_al_u2647_o}),
    .c({_al_u3835_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3836_o,_al_u3835_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*~A)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~C*B*~A)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3838|_al_u3837  (
    .a({open_n29403,_al_u1643_o}),
    .b({open_n29404,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u3837_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u3838_o,_al_u3837_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+~(D)*B*~(C)+D*B*~(C)+~(D)*~(B)*C+~(D)*B*C)"),
    //.LUTF1("(C*A*~(D*B))"),
    //.LUTG0("(D*~(B)*~(C)+~(D)*B*~(C)+D*B*~(C)+~(D)*~(B)*C+~(D)*B*C)"),
    //.LUTG1("(C*A*~(D*B))"),
    .INIT_LUTF0(16'b0000111111111100),
    .INIT_LUTF1(16'b0010000010100000),
    .INIT_LUTG0(16'b0000111111111100),
    .INIT_LUTG1(16'b0010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3840|_al_u3839  (
    .a({_al_u3839_o,open_n29429}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({_al_u2868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,_al_u2767_o}),
    .f({_al_u3840_o,_al_u3839_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(B*~(C@D))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(B*~(C@D))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000001100),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3841|_al_u3842  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,_al_u3841_o}),
    .f({_al_u3841_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~D*~(C*B)))"),
    //.LUT1("(~D*~(~A*~(~C*~B)))"),
    .INIT_LUT0(16'b0101010101000000),
    .INIT_LUT1(16'b0000000010101011),
    .MODE("LOGIC"))
    \_al_u3845|_al_u3844  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm6ow6_lutinv ,_al_u2369_o}),
    .b({_al_u3844_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3845_o,_al_u3844_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(~(A)*~(B)*~(D)+A*~(B)*~(D)+~(A)*B*D))"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("(C*(~(A)*~(B)*~(D)+A*~(B)*~(D)+~(A)*B*D))"),
    //.LUTG1("(~A*~(D*C*B))"),
    .INIT_LUTF0(16'b0100000000110000),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b0100000000110000),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3847|_al_u3846  (
    .a({_al_u3846_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3847_o,_al_u3846_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(A*~(~C*~B)))"),
    //.LUTF1("(~B*A*~(D*~C))"),
    //.LUTG0("(~D*~(A*~(~C*~B)))"),
    //.LUTG1("(~B*A*~(D*~C))"),
    .INIT_LUTF0(16'b0000000001010111),
    .INIT_LUTF1(16'b0010000000100010),
    .INIT_LUTG0(16'b0000000001010111),
    .INIT_LUTG1(16'b0010000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3848|_al_u3849  (
    .a({_al_u3843_o,_al_u3836_o}),
    .b({_al_u3845_o,_al_u3838_o}),
    .c({_al_u3847_o,_al_u3848_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u3848_o,_al_u3849_o}));
  // ../RTL/cortexm0ds_logic.v(18708)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(~D*(C@B)))"),
    //.LUT1("(~B*(A*~(C)*~(D)+~(A)*C*~(D)+A*C*~(D)+A*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010101111101),
    .INIT_LUT1(16'b0010000000110010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3851|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 ,_al_u3309_o}),
    .b({_al_u2790_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zbjiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ncjiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gcjiu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u3314_o,_al_u2790_o}),
    .f({_al_u3851_o,open_n29561}),
    .q({open_n29565,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }));  // ../RTL/cortexm0ds_logic.v(18708)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~D*(C@B))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000000111100),
    .MODE("LOGIC"))
    \_al_u3853|_al_u3852  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jajiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 }),
    .d({_al_u2783_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 }),
    .f({_al_u3853_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jajiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0011000000111111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0011000000111111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3856|_al_u3855  (
    .a({_al_u3854_o,open_n29588}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 ,_al_u1803_o}),
    .c({_al_u3855_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u3856_o,_al_u3855_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u3857|_al_u3557  (
    .a({_al_u3853_o,open_n29613}),
    .b({_al_u3856_o,open_n29614}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot7ow6 }),
    .f({_al_u3857_o,_al_u3557_o}));
  // ../RTL/cortexm0ds_logic.v(17286)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(~B*A*~(D*~C))"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(~B*A*~(D*~C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b0010000000100010),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b0010000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3859|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6_reg  (
    .a({_al_u3857_o,open_n29635}),
    .b({_al_u3858_o,open_n29636}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yb8iu6 ,_al_u3859_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F58iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 ,_al_u3851_o}),
    .f({_al_u3859_o,open_n29654}),
    .q({open_n29658,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 }));  // ../RTL/cortexm0ds_logic.v(17286)
  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u385|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b7  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in }),
    .mi({open_n29666,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 ,_al_u388_o}),
    .q({open_n29681,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [7]}));  // ../RTL/cmsdk_apb_uart.v(603)
  // ../RTL/cortexm0ds_logic.v(18823)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3861|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1qax6_reg  (
    .c({_al_u3603_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u3601_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv }),
    .mi({open_n29696,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 }),
    .q({open_n29701,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] }));  // ../RTL/cortexm0ds_logic.v(18823)
  // ../RTL/cortexm0ds_logic.v(20251)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*D))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("~(~C*~(B*D))"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011110000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1111110011110000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3874|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rekbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 ,open_n29702}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 }),
    .c({_al_u1299_o,\u_cmsdk_mcu/SYSRESETREQ }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9qow6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3874_o,open_n29720}),
    .q({open_n29724,\u_cmsdk_mcu/SYSRESETREQ }));  // ../RTL/cortexm0ds_logic.v(20251)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3877|_al_u3878  (
    .b({_al_u2832_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfiiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aaiiu6 ,_al_u2827_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfiiu6 ,_al_u3878_o}));
  // ../RTL/cortexm0ds_logic.v(18703)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011100100010),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1111011100100010),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3879|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6_reg  (
    .a({open_n29751,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D8iiu6 }),
    .b({_al_u2841_o,_al_u3879_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ,_al_u3880_o}),
    .clk(XTAL1_wire),
    .d({_al_u3878_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 }),
    .f({_al_u3879_o,open_n29770}),
    .q({open_n29774,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 }));  // ../RTL/cortexm0ds_logic.v(18703)
  // ../RTL/cmsdk_apb_uart.v(614)
  EG_PHY_MSLICE #(
    //.LUT0("(D*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u387|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0],open_n29775}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [1]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_in }),
    .q({open_n29791,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [6]}));  // ../RTL/cmsdk_apb_uart.v(614)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u3880|_al_u2920  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 ,open_n29794}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lgkax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkax6 }),
    .d({_al_u3423_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf7ju6 }),
    .f({_al_u3880_o,_al_u2920_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u3885|_al_u3884  (
    .a({open_n29815,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1533_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30],_al_u3797_o}),
    .d({_al_u3884_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [28]}),
    .f({_al_u3885_o,_al_u3884_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3887|_al_u3886  (
    .a({open_n29836,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [30]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/If3pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32]}),
    .f({_al_u3887_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/If3pw6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u3889|_al_u3888  (
    .a({open_n29861,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1541_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [29]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd4pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31]}),
    .f({_al_u3889_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd4pw6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~D*C*A))"),
    //.LUT1("(~C*~(~A*~(~D*B)))"),
    .INIT_LUT0(16'b0011001100010011),
    .INIT_LUT1(16'b0000101000001110),
    .MODE("LOGIC"))
    \_al_u3893|_al_u3892  (
    .a({_al_u3891_o,_al_u696_o}),
    .b({_al_u681_o,_al_u909_o}),
    .c({_al_u3892_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u3893_o,_al_u3892_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~C*~A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(D*~C*~A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011001000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011001000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3895|_al_u3897  (
    .a({open_n29902,_al_u3895_o}),
    .b({_al_u2832_o,_al_u3896_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,_al_u1812_o}),
    .d({_al_u2771_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3895_o,_al_u3897_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3896|_al_u1666  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv }),
    .f({_al_u3896_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vs0iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u3898|_al_u3016  (
    .a({_al_u1269_o,open_n29953}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ,open_n29954}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u3898_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("~(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("~(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0001101110111011),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0001101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3899|_al_u3634  (
    .a({_al_u3109_o,open_n29975}),
    .b({_al_u3898_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv }),
    .c({_al_u2779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv ,_al_u696_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fy8ow6_lutinv ,_al_u3634_o}));
  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u389|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b0  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .clk(XTAL1_wire),
    .d({_al_u388_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ,open_n30020}),
    .q({open_n30024,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [0]}));  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(D*C))"),
    //.LUTF1("(C*A*~(~D*~B))"),
    //.LUTG0("(~B*~A*~(D*C))"),
    //.LUTG1("(C*A*~(~D*~B))"),
    .INIT_LUTF0(16'b0000000100010001),
    .INIT_LUTF1(16'b1010000010000000),
    .INIT_LUTG0(16'b0000000100010001),
    .INIT_LUTG1(16'b1010000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3900|_al_u3894  (
    .a({_al_u3894_o,_al_u2846_o}),
    .b({_al_u3897_o,_al_u3893_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fy8ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8oiu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u3900_o,_al_u3894_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*~A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3901|_al_u3904  (
    .a({open_n30049,_al_u3901_o}),
    .b({open_n30050,_al_u3903_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({_al_u2371_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3901_o,_al_u3904_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*~C))"),
    //.LUT1("(~A*~(~D*~C*B))"),
    .INIT_LUT0(16'b0100010001000000),
    .INIT_LUT1(16'b0101010101010001),
    .MODE("LOGIC"))
    \_al_u3903|_al_u3902  (
    .a({_al_u3902_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3903_o,_al_u3902_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(~D*C))"),
    //.LUT1("(D*C*~(~B*A))"),
    .INIT_LUT0(16'b1000100000001000),
    .INIT_LUT1(16'b1101000000000000),
    .MODE("LOGIC"))
    \_al_u3906|_al_u3905  (
    .a({_al_u3904_o,_al_u2369_o}),
    .b({_al_u3905_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({_al_u2364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u3906_o,_al_u3905_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000011101010),
    .MODE("LOGIC"))
    \_al_u3907|_al_u4001  (
    .a({_al_u3906_o,open_n30111}),
    .b({_al_u2373_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 }),
    .c({_al_u3831_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ,_al_u2373_o}),
    .f({_al_u3907_o,_al_u4001_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u3909|_al_u3908  (
    .a({_al_u3908_o,open_n30132}),
    .b({_al_u2367_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 }),
    .f({_al_u3909_o,_al_u3908_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~B*A*~(D*C))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"))
    \_al_u3911|_al_u3910  (
    .a({_al_u3909_o,_al_u2364_o}),
    .b({_al_u3910_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({_al_u2373_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3911_o,_al_u3910_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3913|_al_u3912  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u3912_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yj8ow6 ,_al_u3912_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D)"),
    //.LUT1("(A*~(C*~(~D*B)))"),
    .INIT_LUT0(16'b0000001101011111),
    .INIT_LUT1(16'b0000101010001010),
    .MODE("LOGIC"))
    \_al_u3915|_al_u3914  (
    .a({_al_u3911_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yj8ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({_al_u3914_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u3915_o,_al_u3914_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~(B*~A))"),
    //.LUT1("(~D*~C*~(B*~A))"),
    .INIT_LUT0(16'b0000000000001011),
    .INIT_LUT1(16'b0000000000001011),
    .MODE("LOGIC"))
    \_al_u3916|_al_u3921  (
    .a({_al_u3907_o,_al_u3916_o}),
    .b({_al_u3915_o,_al_u3920_o}),
    .c({_al_u1812_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u3916_o,_al_u3921_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~B*~(~D*C)))"),
    //.LUTF1("(~D*~C*B*~A)"),
    //.LUTG0("(A*~(~B*~(~D*C)))"),
    //.LUTG1("(~D*~C*B*~A)"),
    .INIT_LUTF0(16'b1000100010101000),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b1000100010101000),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3920|_al_u3919  (
    .a({_al_u3827_o,_al_u1806_o}),
    .b({_al_u3918_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ly2ju6 }),
    .c({_al_u697_o,_al_u604_o}),
    .d({_al_u3919_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u3920_o,_al_u3919_o}));
  // ../RTL/cortexm0ds_logic.v(17735)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*~(~D*~A))"),
    //.LUT1("(D*~(~A*~(C*~B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111101),
    .INIT_LUT1(16'b1011101000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3922|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u3900_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,_al_u3921_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,_al_u3922_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3922_o,open_n30276}),
    .q({open_n30280,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }));  // ../RTL/cortexm0ds_logic.v(17735)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u3925|_al_u3924  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 ,open_n30283}),
    .c({_al_u3924_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u1346_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u3925_o,_al_u3924_o}));
  // ../RTL/cortexm0ds_logic.v(17193)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(B*~(~D*~(C*A)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(B*~(~D*~(C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1100110010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1100110010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3927|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6_reg  (
    .a({_al_u1777_o,open_n30304}),
    .b({_al_u3926_o,_al_u3518_o}),
    .c({_al_u3520_o,_al_u3927_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3927_o,open_n30322}),
    .q({open_n30326,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaipw6 }));  // ../RTL/cortexm0ds_logic.v(17193)
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*A))"),
    //.LUTF1("(B*~(~D*~(C*A)))"),
    //.LUTG0("(~(~D*C)*~(B*A))"),
    //.LUTG1("(B*~(~D*~(C*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011100000111),
    .INIT_LUTF1(16'b1100110010000000),
    .INIT_LUTG0(16'b0111011100000111),
    .INIT_LUTG1(16'b1100110010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3932|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b1  (
    .a({_al_u1777_o,\u_cmsdk_mcu/HWDATA [1]}),
    .b({_al_u3931_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 }),
    .mi({open_n30330,\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3932_o,_al_u3456_o}),
    .q({open_n30345,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [1]}));  // ../RTL/gpio_apbif.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~(C*B)))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(A*~(~D*~(C*B)))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b1010101010000000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1010101010000000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3934|_al_u3935  (
    .a({open_n30346,_al_u3934_o}),
    .b({_al_u3337_o,_al_u1777_o}),
    .c({_al_u3925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 }),
    .f({_al_u3934_o,_al_u3935_o}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(D*A))"),
    //.LUT1("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000011000000),
    .INIT_LUT1(16'b0011111100001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3937|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b10  (
    .a({_al_u1777_o,\u_cmsdk_mcu/HWDATA [10]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcgiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [10]}),
    .c({_al_u3925_o,_al_u3937_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .mi({open_n30381,\u_cmsdk_mcu/HWDATA [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3937_o,_al_u3938_o}),
    .q({open_n30385,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [10]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~(D*A))"),
    //.LUTF1("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("(C*~B*~(D*A))"),
    //.LUTG1("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000000110000),
    .INIT_LUTF1(16'b0011111100001000),
    .INIT_LUTG0(16'b0001000000110000),
    .INIT_LUTG1(16'b0011111100001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3940|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b12  (
    .a({_al_u1777_o,\u_cmsdk_mcu/HWDATA [12]}),
    .b({_al_u3443_o,_al_u3440_o}),
    .c({_al_u3925_o,_al_u3940_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W51bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .mi({open_n30389,\u_cmsdk_mcu/HWDATA [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3940_o,_al_u3941_o}),
    .q({open_n30404,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [12]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cortexm0ds_logic.v(19455)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(A*~(~D*~(C*B)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1010101010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1010101010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3944|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6_reg  (
    .a({_al_u3943_o,open_n30405}),
    .b({_al_u1777_o,_al_u3492_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzfiu6_lutinv ,_al_u3944_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3944_o,open_n30423}),
    .q({open_n30427,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/At2bx6 }));  // ../RTL/cortexm0ds_logic.v(19455)
  // ../RTL/cortexm0ds_logic.v(19431)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1010101010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3947|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6_reg  (
    .a({_al_u3946_o,open_n30428}),
    .b({_al_u1777_o,_al_u3498_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mxfiu6_lutinv ,_al_u3947_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3947_o,open_n30442}),
    .q({open_n30446,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok2bx6 }));  // ../RTL/cortexm0ds_logic.v(19431)
  // ../RTL/cortexm0ds_logic.v(19467)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1010101010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3950|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6_reg  (
    .a({_al_u3949_o,open_n30447}),
    .b({_al_u1777_o,_al_u3503_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivfiu6_lutinv ,_al_u3950_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3950_o,open_n30461}),
    .q({open_n30465,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx2bx6 }));  // ../RTL/cortexm0ds_logic.v(19467)
  // ../RTL/cortexm0ds_logic.v(19479)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(A*~(~D*~(C*B)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1010101010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1010101010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3953|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6_reg  (
    .a({_al_u3952_o,open_n30466}),
    .b({_al_u1777_o,_al_u3508_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv ,_al_u3953_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3953_o,open_n30484}),
    .q({open_n30488,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M13bx6 }));  // ../RTL/cortexm0ds_logic.v(19479)
  // ../RTL/cortexm0ds_logic.v(19491)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(B*~(~D*~(C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1100110010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3956|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6_reg  (
    .a({_al_u1777_o,open_n30489}),
    .b({_al_u3955_o,_al_u3513_o}),
    .c({_al_u3515_o,_al_u3956_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3956_o,open_n30503}),
    .q({open_n30507,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S53bx6 }));  // ../RTL/cortexm0ds_logic.v(19491)
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~C)*~(B*A))"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111011101110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3958|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b6  (
    .a({open_n30508,\u_cmsdk_mcu/HWDATA [6]}),
    .b({_al_u3359_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({_al_u3925_o,_al_u3359_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 }),
    .mi({open_n30519,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3958_o,_al_u3360_o}),
    .q({open_n30523,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6]}));  // ../RTL/gpio_apbif.v(303)
  // ../RTL/cortexm0ds_logic.v(19824)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*B))"),
    //.LUT1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000001010000),
    .INIT_LUT1(16'b1010101010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3959|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6_reg  (
    .a({_al_u3958_o,_al_u3874_o}),
    .b({_al_u1777_o,\u_cmsdk_mcu/HWDATA [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv ,_al_u3959_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3959_o,open_n30537}),
    .q({open_n30541,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp9bx6 }));  // ../RTL/cortexm0ds_logic.v(19824)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u395|_al_u6302  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ,_al_u6302_o}));
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~C)*~(B*A))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~(~D*~C)*~(B*A))"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011101110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0111011101110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3961|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b7  (
    .a({open_n30570,\u_cmsdk_mcu/HWDATA [7]}),
    .b({_al_u3369_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({_al_u3925_o,_al_u3369_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({_al_u3372_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 }),
    .mi({open_n30574,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3961_o,_al_u3370_o}),
    .q({open_n30589,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7]}));  // ../RTL/gpio_apbif.v(303)
  // ../RTL/cortexm0ds_logic.v(19539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*B))"),
    //.LUT1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000001010000),
    .INIT_LUT1(16'b1010101010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3962|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6_reg  (
    .a({_al_u3961_o,_al_u3874_o}),
    .b({_al_u1777_o,\u_cmsdk_mcu/HWDATA [7]}),
    .c({_al_u3372_o,_al_u3962_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3962_o,open_n30603}),
    .q({open_n30607,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Om3bx6 }));  // ../RTL/cortexm0ds_logic.v(19539)
  // ../RTL/cortexm0ds_logic.v(19347)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~A)"),
    //.LUTF1("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("(D*~C*~B*~A)"),
    //.LUTG1("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0011111100001000),
    .INIT_LUTG0(16'b0000000100000000),
    .INIT_LUTG1(16'b0011111100001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3964|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6_reg  (
    .a({_al_u1777_o,_al_u3874_o}),
    .b({_al_u3454_o,_al_u3449_o}),
    .c({_al_u3925_o,_al_u3450_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 ,_al_u3964_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3964_o,open_n30625}),
    .q({open_n30629,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1bx6 }));  // ../RTL/cortexm0ds_logic.v(19347)
  // ../RTL/cortexm0ds_logic.v(19371)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1010101010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3967|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6_reg  (
    .a({_al_u3966_o,open_n30630}),
    .b({_al_u1777_o,_al_u3461_o}),
    .c({_al_u3463_o,_al_u3967_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3967_o,open_n30644}),
    .q({open_n30648,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz1bx6 }));  // ../RTL/cortexm0ds_logic.v(19371)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3969|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b3  (
    .b({_al_u3925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n277 ),
    .clk(XTAL1_wire),
    .d({_al_u3468_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3969_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [3]}),
    .q({open_n30666,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u396|_al_u550  (
    .a({open_n30667,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 }));
  // ../RTL/cortexm0ds_logic.v(19383)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(A*~(~D*~(C*B)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1010101010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1010101010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3970|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6_reg  (
    .a({_al_u3969_o,open_n30688}),
    .b({_al_u1777_o,_al_u3466_o}),
    .c({_al_u3468_o,_al_u3970_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3970_o,open_n30706}),
    .q({open_n30710,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S32bx6 }));  // ../RTL/cortexm0ds_logic.v(19383)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3972|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b4  (
    .b({_al_u3925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [4]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n279 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3972_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [4]}),
    .q({open_n30728,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cortexm0ds_logic.v(19407)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(A*~(~D*~(C*B)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1010101010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1010101010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3973|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6_reg  (
    .a({_al_u3972_o,open_n30729}),
    .b({_al_u1777_o,_al_u3471_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhdiu6_lutinv ,_al_u3973_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3973_o,open_n30747}),
    .q({open_n30751,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cc2bx6 }));  // ../RTL/cortexm0ds_logic.v(19407)
  // ../RTL/cortexm0ds_logic.v(19419)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(A*~(~D*~(C*B)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1010101010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1010101010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3976|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6_reg  (
    .a({_al_u3975_o,open_n30752}),
    .b({_al_u1777_o,_al_u3477_o}),
    .c({_al_u3479_o,_al_u3976_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3976_o,open_n30770}),
    .q({open_n30774,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ig2bx6 }));  // ../RTL/cortexm0ds_logic.v(19419)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3978|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg7_b6  (
    .b({_al_u3925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n283 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3978_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [6]}),
    .q({open_n30796,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6]}));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cortexm0ds_logic.v(20025)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(A*~(~D*~(C*B)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1010101010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1010101010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3979|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6_reg  (
    .a({_al_u3978_o,open_n30797}),
    .b({_al_u1777_o,_al_u3482_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv ,_al_u3979_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3979_o,open_n30815}),
    .q({open_n30819,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vyfbx6 }));  // ../RTL/cortexm0ds_logic.v(20025)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u397|_al_u1303  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }));
  // ../RTL/cortexm0ds_logic.v(19443)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1010101010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3982|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6_reg  (
    .a({_al_u3981_o,open_n30848}),
    .b({_al_u1777_o,_al_u3487_o}),
    .c({_al_u3489_o,_al_u3982_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3982_o,open_n30862}),
    .q({open_n30866,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uo2bx6 }));  // ../RTL/cortexm0ds_logic.v(19443)
  // ../RTL/cortexm0ds_logic.v(19503)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(B*~(~D*~(C*A)))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(B*~(~D*~(C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b1100110010000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b1100110010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3985|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6_reg  (
    .a({_al_u1777_o,open_n30867}),
    .b({_al_u3984_o,_al_u3528_o}),
    .c({_al_u3530_o,_al_u3985_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3985_o,open_n30885}),
    .q({open_n30889,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y93bx6 }));  // ../RTL/cortexm0ds_logic.v(19503)
  // ../RTL/cortexm0ds_logic.v(19515)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(B*~(~D*~(C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1100110010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3988|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6_reg  (
    .a({_al_u1777_o,open_n30890}),
    .b({_al_u3987_o,_al_u3523_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 ,_al_u3988_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 ,_al_u3874_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3988_o,open_n30904}),
    .q({open_n30908,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ee3bx6 }));  // ../RTL/cortexm0ds_logic.v(19515)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(C*~(B*D))"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3990|_al_u574  (
    .a({open_n30909,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [1]}),
    .b({_al_u3925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .d({_al_u3335_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .f({_al_u3990_o,_al_u574_o}));
  // ../RTL/cortexm0ds_logic.v(19275)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(D*B))"),
    //.LUTF1("(A*~(~D*~(C*B)))"),
    //.LUTG0("(C*~A*~(D*B))"),
    //.LUTG1("(A*~(~D*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000001010000),
    .INIT_LUTF1(16'b1010101010000000),
    .INIT_LUTG0(16'b0001000001010000),
    .INIT_LUTG1(16'b1010101010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3991|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6_reg  (
    .a({_al_u3990_o,_al_u3874_o}),
    .b({_al_u1777_o,\u_cmsdk_mcu/HWDATA [0]}),
    .c({_al_u3335_o,_al_u3991_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3991_o,open_n30951}),
    .q({open_n30955,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S11bx6 }));  // ../RTL/cortexm0ds_logic.v(19275)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3994|_al_u3993  (
    .b({open_n30958,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u3993_o,_al_u909_o}),
    .f({_al_u3994_o,_al_u3993_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~D*~B*~(C*A))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000000010011),
    .MODE("LOGIC"))
    \_al_u3996|_al_u3995  (
    .a({_al_u3183_o,open_n30983}),
    .b({_al_u3994_o,_al_u1582_o}),
    .c({_al_u3910_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u3995_o,_al_u679_o}),
    .f({_al_u3996_o,_al_u3995_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3998|_al_u3997  (
    .b({_al_u3997_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8ziu6 ,_al_u3997_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D*A)))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .INIT_LUT0(16'b0010001100000011),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"))
    \_al_u4000|_al_u3999  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dd7ow6 ,_al_u2371_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8ziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({_al_u3246_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ea7ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .f({_al_u4000_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ea7ow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~C*A*~(~D*~B))"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000101000001000),
    .MODE("LOGIC"))
    \_al_u4003|_al_u4002  (
    .a({_al_u3996_o,_al_u1812_o}),
    .b({_al_u4000_o,_al_u4001_o}),
    .c({_al_u4002_o,_al_u2369_o}),
    .d({_al_u1812_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u4003_o,_al_u4002_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~C*B))"),
    //.LUT1("(A*~(D*C*~B))"),
    .INIT_LUT0(16'b1010001010101010),
    .INIT_LUT1(16'b1000101010101010),
    .MODE("LOGIC"))
    \_al_u4004|_al_u4413  (
    .a({_al_u4003_o,_al_u4412_o}),
    .b({_al_u3109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .c({_al_u1806_o,_al_u3109_o}),
    .d({_al_u1266_o,_al_u1266_o}),
    .f({_al_u4004_o,_al_u4413_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(~(B)*~(C)*~(D)+~(B)*C*~(D)+B*C*~(D)+B*~(C)*D+B*C*D))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1000100010100010),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u4005|_al_u4375  (
    .a({open_n31086,_al_u4374_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbkiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .d({_al_u3227_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh7ow6 ,_al_u4375_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~(B*~A))"),
    //.LUTF1("(~D*~(C*~B*A))"),
    //.LUTG0("(~D*~C*~(B*~A))"),
    //.LUTG1("(~D*~(C*~B*A))"),
    .INIT_LUTF0(16'b0000000000001011),
    .INIT_LUTF1(16'b0000000011011111),
    .INIT_LUTG0(16'b0000000000001011),
    .INIT_LUTG1(16'b0000000011011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4009|_al_u4008  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qz0ju6 ,_al_u4007_o}),
    .b({_al_u4008_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u4009_o,_al_u4008_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(A*~(C*~(~D*~B)))"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b0000101000101010),
    .MODE("LOGIC"))
    \_al_u4010|_al_u4006  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yd7ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh7ow6 }),
    .b({_al_u4009_o,_al_u4001_o}),
    .c({_al_u2365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmiiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u4010_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yd7ow6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17623)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*~A))"),
    //.LUTF1("(~D*~(A*~(C*~B)))"),
    //.LUTG0("(~(~D*C)*~(B*~A))"),
    //.LUTG1("(~D*~(A*~(C*~B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b0000000001110101),
    .INIT_LUTG0(16'b1011101100001011),
    .INIT_LUTG1(16'b0000000001110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4011|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6_reg  (
    .a({_al_u4004_o,_al_u4011_o}),
    .b({_al_u4010_o,_al_u4023_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uyiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4011_o,open_n31168}),
    .q({open_n31172,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }));  // ../RTL/cortexm0ds_logic.v(17623)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~B*~(~D*~C)))"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1000100010001010),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u4012|_al_u2646  (
    .a({open_n31173,_al_u1658_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4012_o,_al_u2646_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~A*~(D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~A*~(D*B))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000100000101),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4013|_al_u3657  (
    .a({_al_u3189_o,open_n31194}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv ,open_n31195}),
    .c({_al_u4012_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({_al_u1582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv }),
    .f({_al_u4013_o,_al_u3657_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4014|_al_u2392  (
    .a({_al_u904_o,open_n31220}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,open_n31221}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u2392_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u4014_o,_al_u2392_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*C*~B*A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u4015|_al_u3656  (
    .a({_al_u4013_o,open_n31246}),
    .b({_al_u3186_o,open_n31247}),
    .c({_al_u4014_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu9ow6_lutinv ,_al_u1346_o}),
    .f({_al_u4015_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(~D*~C*~B*A)"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"))
    \_al_u4018|_al_u4016  (
    .a({_al_u4015_o,open_n31268}),
    .b({_al_u1784_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u4016_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u4017_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu9ow6 }),
    .f({_al_u4018_o,_al_u4016_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4019|_al_u1268  (
    .b({_al_u1268_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u1802_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us2ju6 }),
    .f({_al_u4019_o,_al_u1268_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u401|_al_u4047  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5eiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~A)"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(D*~C*~B*~A)"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0000000100000000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4021|_al_u4020  (
    .a({_al_u4018_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .b({_al_u4019_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V17ow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u4021_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V17ow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"))
    \_al_u4022|_al_u908  (
    .a({_al_u908_o,open_n31367}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ,open_n31368}),
    .c({_al_u932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv }),
    .f({_al_u4022_o,_al_u908_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(A*~(~D*~(C*~B)))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1010101000100000),
    .MODE("LOGIC"))
    \_al_u4023|_al_u3824  (
    .a({_al_u4021_o,open_n31389}),
    .b({_al_u3824_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .c({_al_u4022_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv }),
    .f({_al_u4023_o,_al_u3824_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4026|_al_u4239  (
    .b({open_n31412,_al_u1250_o}),
    .c({_al_u4025_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 ,_al_u4239_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~(~D*~A))"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(~C*B*~(~D*~A))"),
    //.LUTG1("(C*~(B*D))"),
    .INIT_LUTF0(16'b0000110000001000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b0000110000001000),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4028|_al_u2306  (
    .a({open_n31433,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 }),
    .b({_al_u4027_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6yhu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,_al_u2305_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .f({_al_u4028_o,_al_u2306_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4029|_al_u1253  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ,open_n31458}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 }),
    .f({_al_u4029_o,_al_u1253_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .INIT_LUTF0(16'b0001101111110000),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b0001101111110000),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4031|_al_u4030  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .b({_al_u4029_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .c({_al_u4030_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }),
    .f({_al_u4031_o,_al_u4030_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~B*(D@A)))"),
    //.LUT1("(D*~(C*~B*~A))"),
    .INIT_LUT0(16'b0000111000001101),
    .INIT_LUT1(16'b1110111100000000),
    .MODE("LOGIC"))
    \_al_u4032|_al_u3430  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbyhu6 ,_al_u1756_o}),
    .b({_al_u4028_o,_al_u1761_o}),
    .c({_al_u4031_o,_al_u1763_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .f({_al_u4032_o,_al_u3430_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4035|_al_u4034  (
    .a({open_n31527,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1397_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13],_al_u3797_o}),
    .d({_al_u4034_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [11]}),
    .f({_al_u4035_o,_al_u4034_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*A*~(~D*~C))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0010001000100000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u4039|_al_u4038  (
    .a({_al_u4037_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zyoiu6 }),
    .b({_al_u4038_o,_al_u1812_o}),
    .c({_al_u697_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u3667_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u4039_o,_al_u4038_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~D*~(B*~A)))"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(~C*~(~D*~(B*~A)))"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b0000111100000100),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000111100000100),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4040|_al_u4049  (
    .a({open_n31572,_al_u4040_o}),
    .b({_al_u4039_o,_al_u4046_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,_al_u4048_o}),
    .d({_al_u4036_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({_al_u4040_o,_al_u4049_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u4043|_al_u4041  (
    .a({_al_u4041_o,open_n31597}),
    .b({_al_u4042_o,_al_u604_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u3110_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .f({_al_u4043_o,_al_u4041_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*A*~(~D*B))"),
    //.LUT1("(D*C*~(~B*A))"),
    .INIT_LUT0(16'b0000101000000010),
    .INIT_LUT1(16'b1101000000000000),
    .MODE("LOGIC"))
    \_al_u4045|_al_u4046  (
    .a({_al_u1812_o,_al_u4043_o}),
    .b({_al_u4044_o,_al_u2754_o}),
    .c({_al_u930_o,_al_u4045_o}),
    .d({_al_u1359_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u4045_o,_al_u4046_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*~A*~(~D*B))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*~A*~(~D*B))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0101000000010000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0101000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4050|_al_u2860  (
    .a({_al_u4049_o,open_n31638}),
    .b({_al_u2860_o,open_n31639}),
    .c({_al_u903_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u3811_o,_al_u1812_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,_al_u2860_o}));
  // ../RTL/cortexm0ds_logic.v(18276)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4052|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6_reg  (
    .a({open_n31664,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emmiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 }),
    .mi({open_n31668,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .f({_al_u4052_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emmiu6 }),
    .q({open_n31684,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 }));  // ../RTL/cortexm0ds_logic.v(18276)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4056|_al_u4055  (
    .a({open_n31685,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1429_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17],_al_u3797_o}),
    .d({_al_u4055_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [15]}),
    .f({_al_u4056_o,_al_u4055_o}));
  // ../RTL/cortexm0ds_logic.v(17814)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4058|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbmiu6 ,_al_u4058_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,_al_u4056_o}),
    .f({_al_u4058_o,open_n31722}),
    .q({open_n31726,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 }));  // ../RTL/cortexm0ds_logic.v(17814)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u405|_al_u3266  (
    .b({open_n31729,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 }),
    .f({_al_u405_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4061|_al_u4060  (
    .a({open_n31750,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1437_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18],_al_u3797_o}),
    .d({_al_u4060_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [16]}),
    .f({_al_u4061_o,_al_u4060_o}));
  // ../RTL/cortexm0ds_logic.v(19937)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4063|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6_reg  (
    .a({open_n31771,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8miu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 }),
    .mi({open_n31782,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .f({_al_u4063_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8miu6 }),
    .q({open_n31787,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 }));  // ../RTL/cortexm0ds_logic.v(19937)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4066|_al_u4065  (
    .a({open_n31788,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1445_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19],_al_u3797_o}),
    .d({_al_u4065_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [17]}),
    .f({_al_u4066_o,_al_u4065_o}));
  // ../RTL/cortexm0ds_logic.v(18316)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4068|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6_reg  (
    .a({open_n31813,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5miu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 }),
    .mi({open_n31824,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 }),
    .f({_al_u4068_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5miu6 }),
    .q({open_n31829,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 }));  // ../RTL/cortexm0ds_logic.v(18316)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4071|_al_u4070  (
    .a({open_n31830,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1453_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20],_al_u3797_o}),
    .d({_al_u4070_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [18]}),
    .f({_al_u4071_o,_al_u4070_o}));
  // ../RTL/cortexm0ds_logic.v(18249)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4073|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6_reg  (
    .a({open_n31855,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2miu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 }),
    .mi({open_n31866,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .f({_al_u4073_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2miu6 }),
    .q({open_n31871,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 }));  // ../RTL/cortexm0ds_logic.v(18249)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4076|_al_u4075  (
    .a({open_n31872,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1461_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21],_al_u3797_o}),
    .d({_al_u4075_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [19]}),
    .f({_al_u4076_o,_al_u4075_o}));
  // ../RTL/cortexm0ds_logic.v(19978)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4078|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6_reg  (
    .a({open_n31893,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hzliu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 }),
    .mi({open_n31904,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .f({_al_u4078_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hzliu6 }),
    .q({open_n31909,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 }));  // ../RTL/cortexm0ds_logic.v(19978)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4081|_al_u4080  (
    .a({open_n31910,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1469_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22],_al_u3797_o}),
    .d({_al_u4080_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [20]}),
    .f({_al_u4081_o,_al_u4080_o}));
  // ../RTL/cortexm0ds_logic.v(19990)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4083|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6_reg  (
    .a({open_n31931,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwliu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 }),
    .mi({open_n31935,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .f({_al_u4083_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwliu6 }),
    .q({open_n31951,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 }));  // ../RTL/cortexm0ds_logic.v(19990)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4086|_al_u4085  (
    .a({open_n31952,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1477_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23],_al_u3797_o}),
    .d({_al_u4085_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [21]}),
    .f({_al_u4086_o,_al_u4085_o}));
  // ../RTL/cortexm0ds_logic.v(19996)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4088|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctliu6 ,_al_u4088_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,_al_u4086_o}),
    .f({_al_u4088_o,open_n31993}),
    .q({open_n31997,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 }));  // ../RTL/cortexm0ds_logic.v(19996)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u408|_al_u5001  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjyiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ,_al_u5001_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4091|_al_u4090  (
    .a({open_n32026,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1485_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24],_al_u3797_o}),
    .d({_al_u4090_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [22]}),
    .f({_al_u4091_o,_al_u4090_o}));
  // ../RTL/cortexm0ds_logic.v(20102)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4093|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6_reg  (
    .a({open_n32051,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kv9iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 }),
    .mi({open_n32062,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .f({_al_u4093_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kv9iu6 }),
    .q({open_n32067,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 }));  // ../RTL/cortexm0ds_logic.v(20102)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(~B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000110111011101),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4096|_al_u4095  (
    .a({open_n32068,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27],_al_u3797_o}),
    .d({_al_u4095_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [25]}),
    .f({_al_u4096_o,_al_u4095_o}));
  // ../RTL/cortexm0ds_logic.v(19948)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4098|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6_reg  (
    .a({open_n32089,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzkiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 }),
    .mi({open_n32093,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .f({_al_u4098_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzkiu6 }),
    .q({open_n32109,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 }));  // ../RTL/cortexm0ds_logic.v(19948)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u409|_al_u407  (
    .b({open_n32112,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(~B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000110111011101),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4101|_al_u4100  (
    .a({open_n32137,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28],_al_u3797_o}),
    .d({_al_u4100_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [26]}),
    .f({_al_u4101_o,_al_u4100_o}));
  // ../RTL/cortexm0ds_logic.v(19964)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4103|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6_reg  (
    .a({open_n32158,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2liu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 }),
    .mi({open_n32169,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .f({_al_u4103_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2liu6 }),
    .q({open_n32174,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 }));  // ../RTL/cortexm0ds_logic.v(19964)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4106|_al_u4105  (
    .a({open_n32175,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1608_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9],_al_u3797_o}),
    .d({_al_u4105_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [7]}),
    .f({_al_u4106_o,_al_u4105_o}));
  // ../RTL/cortexm0ds_logic.v(18256)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4108|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6_reg  (
    .a({open_n32200,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3niu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 }),
    .mi({open_n32211,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .f({_al_u4108_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y3niu6 }),
    .q({open_n32216,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 }));  // ../RTL/cortexm0ds_logic.v(18256)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4111|_al_u4110  (
    .a({open_n32217,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1624_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11],_al_u3797_o}),
    .d({_al_u4110_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [9]}),
    .f({_al_u4111_o,_al_u4110_o}));
  // ../RTL/cortexm0ds_logic.v(17855)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4113|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivmiu6 ,_al_u4113_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,_al_u4111_o}),
    .f({_al_u4113_o,open_n32262}),
    .q({open_n32266,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 }));  // ../RTL/cortexm0ds_logic.v(17855)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4116|_al_u4115  (
    .a({open_n32267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1632_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [10]}),
    .d({_al_u4115_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12]}),
    .f({_al_u4116_o,_al_u4115_o}));
  // ../RTL/cortexm0ds_logic.v(19809)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4118|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6_reg  (
    .a({open_n32288,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Womiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 }),
    .mi({open_n32299,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .f({_al_u4118_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Womiu6 }),
    .q({open_n32304,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 }));  // ../RTL/cortexm0ds_logic.v(19809)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u411|_al_u399  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4121|_al_u4120  (
    .a({open_n32329,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1616_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8],_al_u3797_o}),
    .d({_al_u4120_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [6]}),
    .f({_al_u4121_o,_al_u4120_o}));
  // ../RTL/cortexm0ds_logic.v(18171)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4123|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6_reg  (
    .a({open_n32350,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krkiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 }),
    .mi({open_n32354,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 }),
    .f({_al_u4123_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krkiu6 }),
    .q({open_n32370,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 }));  // ../RTL/cortexm0ds_logic.v(18171)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4126|_al_u4125  (
    .a({open_n32371,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1405_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [12]}),
    .d({_al_u4125_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14]}),
    .f({_al_u4126_o,_al_u4125_o}));
  // ../RTL/cortexm0ds_logic.v(18297)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4128|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6_reg  (
    .a({open_n32392,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 }),
    .mi({open_n32403,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .f({_al_u4128_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmiu6 }),
    .q({open_n32408,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 }));  // ../RTL/cortexm0ds_logic.v(18297)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u412|_al_u5031  (
    .b({open_n32411,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ,_al_u5030_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ,_al_u5031_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4131|_al_u4130  (
    .a({open_n32436,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1413_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [13]}),
    .d({_al_u4130_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15]}),
    .f({_al_u4131_o,_al_u4130_o}));
  // ../RTL/cortexm0ds_logic.v(19895)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4133|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6_reg  (
    .a({open_n32461,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ugmiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 }),
    .mi({open_n32465,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .f({_al_u4133_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ugmiu6 }),
    .q({open_n32481,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 }));  // ../RTL/cortexm0ds_logic.v(19895)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4136|_al_u4135  (
    .a({open_n32482,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1421_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [14]}),
    .d({_al_u4135_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16]}),
    .f({_al_u4136_o,_al_u4135_o}));
  // ../RTL/cortexm0ds_logic.v(18296)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4138|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6_reg  (
    .a({open_n32507,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cemiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 }),
    .mi({open_n32511,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .f({_al_u4138_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cemiu6 }),
    .q({open_n32527,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 }));  // ../RTL/cortexm0ds_logic.v(18296)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(~B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000110111011101),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4141|_al_u4140  (
    .a({open_n32528,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7],_al_u3797_o}),
    .d({_al_u4140_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [5]}),
    .f({_al_u4141_o,_al_u4140_o}));
  // ../RTL/cortexm0ds_logic.v(19817)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4143|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6_reg  (
    .a({open_n32549,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zokiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 }),
    .mi({open_n32560,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 }),
    .f({_al_u4143_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zokiu6 }),
    .q({open_n32565,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 }));  // ../RTL/cortexm0ds_logic.v(19817)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u4145|_al_u2812  (
    .b({_al_u2868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 }),
    .f({_al_u4145_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nz2ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*A*~(~C*~B))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*A*~(~C*~B))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1010100000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1010100000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4146|_al_u5854  (
    .a({open_n32588,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .f({_al_u4146_o,_al_u5854_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A*~(~D*B))"),
    //.LUT1("(~B*A*~(D*C))"),
    .INIT_LUT0(16'b0000010100000001),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"))
    \_al_u4147|_al_u5850  (
    .a({_al_u4145_o,_al_u1296_o}),
    .b({_al_u4146_o,_al_u1329_o}),
    .c({_al_u682_o,_al_u1662_o}),
    .d({_al_u1329_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u4147_o,_al_u5850_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(D*~(~C*~B*~A))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(D*~(~C*~B*~A))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111111000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111111000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4148|_al_u694  (
    .a({_al_u604_o,open_n32633}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ,open_n32634}),
    .c({_al_u1336_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u2868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u4148_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u414|_al_u524  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xznow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(A*~(C*~B)))"),
    //.LUT1("(~C*A*~(D*B))"),
    .INIT_LUT0(16'b0000000001110101),
    .INIT_LUT1(16'b0000001000001010),
    .MODE("LOGIC"))
    \_al_u4150|_al_u4149  (
    .a({_al_u4147_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Obbow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u4148_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrcpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u4150_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrcpw6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .INIT_LUTF0(16'b1010001010000000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010001010000000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4152|_al_u4151  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ,_al_u3122_o}),
    .b({_al_u4151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4152_o,_al_u4151_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u4155|_al_u4154  (
    .a({_al_u4150_o,_al_u2849_o}),
    .b({_al_u4152_o,_al_u4153_o}),
    .c({_al_u4154_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({_al_u4155_o,_al_u4154_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~C*~B*~D)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4157|_al_u4156  (
    .a({open_n32747,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .b({_al_u4156_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .d({_al_u1799_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .f({_al_u4157_o,_al_u4156_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*~A)"),
    //.LUT1("(~C*~A*~(D*B))"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0000000100000101),
    .MODE("LOGIC"))
    \_al_u4163|_al_u4162  (
    .a({_al_u4161_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .b({_al_u903_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .c({_al_u4162_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4163_o,_al_u4162_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u4165|_al_u3917  (
    .a({_al_u4163_o,open_n32792}),
    .b({_al_u4164_o,open_n32793}),
    .c({_al_u1269_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({_al_u678_o,_al_u678_o}),
    .f({_al_u4165_o,_al_u3917_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~A*~(~D*B)))"),
    //.LUTF1("(A*~(D*~(C*~B)))"),
    //.LUTG0("(C*~(~A*~(~D*B)))"),
    //.LUTG1("(A*~(D*~(C*~B)))"),
    .INIT_LUTF0(16'b1010000011100000),
    .INIT_LUTF1(16'b0010000010101010),
    .INIT_LUTG0(16'b1010000011100000),
    .INIT_LUTG1(16'b0010000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4166|_al_u4160  (
    .a({_al_u4155_o,_al_u4158_o}),
    .b({_al_u4160_o,_al_u4159_o}),
    .c({_al_u4165_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u4166_o,_al_u4160_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4168|_al_u4289  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u4166_o,_al_u4166_o}),
    .f({_al_u4168_o,_al_u4289_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u416|_al_u548  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u4170|_al_u4169  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 ,_al_u1299_o}),
    .d({_al_u4169_o,_al_u4168_o}),
    .f({_al_u4170_o,_al_u4169_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4173|_al_u4172  (
    .b({open_n32916,_al_u679_o}),
    .c({_al_u4172_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({_al_u4166_o,_al_u3993_o}),
    .f({_al_u4173_o,_al_u4172_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~B*A)"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(D*C*~B*A)"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4176|_al_u4175  (
    .a({open_n32941,_al_u2860_o}),
    .b({_al_u4175_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8fax6 }),
    .d({_al_u4049_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 ,_al_u4175_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*B))"),
    //.LUTF1("(C*~(D*B*A))"),
    //.LUTG0("(~A*~(D*C*B))"),
    //.LUTG1("(C*~(D*B*A))"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b0111000011110000),
    .INIT_LUTG0(16'b0001010101010101),
    .INIT_LUTG1(16'b0111000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4178|_al_u4177  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqoiu6_lutinv ,_al_u2373_o}),
    .b({_al_u1812_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqoiu6 }));
  // ../RTL/cortexm0ds_logic.v(18162)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4181|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6_reg  (
    .a({open_n32990,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwkiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 }),
    .mi({open_n32994,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .f({_al_u4181_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwkiu6 }),
    .q({open_n33010,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 }));  // ../RTL/cortexm0ds_logic.v(18162)
  // ../RTL/cortexm0ds_logic.v(20253)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4182|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6_reg  (
    .b({_al_u4181_o,_al_u4184_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4182_o}),
    .f({_al_u4182_o,open_n33027}),
    .q({open_n33031,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 }));  // ../RTL/cortexm0ds_logic.v(20253)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4184|_al_u4183  (
    .a({open_n33032,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1493_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25],_al_u3797_o}),
    .d({_al_u4183_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [23]}),
    .f({_al_u4184_o,_al_u4183_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u4186|_al_u4179  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpoiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 }));
  // ../RTL/cortexm0ds_logic.v(18161)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4188|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6_reg  (
    .a({open_n33081,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipliu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 }),
    .mi({open_n33092,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .f({_al_u4188_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ipliu6 }),
    .q({open_n33097,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 }));  // ../RTL/cortexm0ds_logic.v(18161)
  // ../RTL/cortexm0ds_logic.v(19940)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4189|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6_reg  (
    .b({_al_u4188_o,_al_u4191_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ,_al_u4189_o}),
    .f({_al_u4189_o,open_n33118}),
    .q({open_n33122,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 }));  // ../RTL/cortexm0ds_logic.v(19940)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u418|_al_u5260  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vynow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ,_al_u5260_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(~B*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*C)*~(~B*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000110111011101),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000110111011101),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4191|_al_u4190  (
    .a({open_n33147,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26],_al_u3797_o}),
    .d({_al_u4190_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [24]}),
    .f({_al_u4191_o,_al_u4190_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u4194|_al_u7168  (
    .a({open_n33172,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocniu6 ,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [27]}),
    .f({_al_u4194_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxbow6 }));
  // ../RTL/cortexm0ds_logic.v(17553)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4195|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6_reg  (
    .b({_al_u4194_o,_al_u4197_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4195_o}),
    .f({_al_u4195_o,open_n33213}),
    .q({open_n33217,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 }));  // ../RTL/cortexm0ds_logic.v(17553)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4197|_al_u4196  (
    .a({open_n33218,_al_u3808_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u1525_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29],_al_u3797_o}),
    .d({_al_u4196_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [27]}),
    .f({_al_u4197_o,_al_u4196_o}));
  // ../RTL/cortexm0ds_logic.v(20106)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4200|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6_reg  (
    .a({open_n33239,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mj8iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 }),
    .mi({open_n33243,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 }),
    .f({_al_u4200_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mj8iu6 }),
    .q({open_n33259,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 }));  // ../RTL/cortexm0ds_logic.v(20106)
  // ../RTL/cortexm0ds_logic.v(18049)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4201|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6_reg  (
    .b({_al_u4200_o,_al_u3885_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4201_o}),
    .f({_al_u4201_o,open_n33276}),
    .q({open_n33280,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 }));  // ../RTL/cortexm0ds_logic.v(18049)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4204|_al_u7165  (
    .a({open_n33281,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8liu6 ,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [29]}),
    .f({_al_u4204_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2cow6 }));
  // ../RTL/cortexm0ds_logic.v(19969)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4205|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6_reg  (
    .b({_al_u4204_o,_al_u3889_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4205_o}),
    .f({_al_u4205_o,open_n33326}),
    .q({open_n33330,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 }));  // ../RTL/cortexm0ds_logic.v(19969)
  // ../RTL/cortexm0ds_logic.v(18404)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4208|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6_reg  (
    .a({open_n33331,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmoiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 }),
    .mi({open_n33335,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .f({_al_u4208_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmoiu6 }),
    .q({open_n33351,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 }));  // ../RTL/cortexm0ds_logic.v(18404)
  // ../RTL/cortexm0ds_logic.v(17477)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4209|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6_reg  (
    .b({_al_u4208_o,_al_u3887_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4209_o}),
    .f({_al_u4209_o,open_n33372}),
    .q({open_n33376,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 }));  // ../RTL/cortexm0ds_logic.v(17477)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u420|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0],_al_u357_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [0],_al_u358_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [0],_al_u359_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [0],_al_u360_o}),
    .mi({open_n33380,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 }),
    .q({open_n33395,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [0]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cortexm0ds_logic.v(18287)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4212|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6_reg  (
    .a({open_n33396,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz8iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B29iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 }),
    .mi({open_n33400,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4212_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz8iu6 }),
    .q({open_n33415,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 }));  // ../RTL/cortexm0ds_logic.v(18287)
  // ../RTL/cortexm0ds_logic.v(20231)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(~A*~(D*~C)))"),
    //.LUTG0("~(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(~A*~(D*~C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110101011000000),
    .INIT_LUTF1(16'b1000110010001000),
    .INIT_LUTG0(16'b1110101011000000),
    .INIT_LUTG1(16'b1000110010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4213|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 ,_al_u3808_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U19iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4213_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 }),
    .q({open_n33435,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 }));  // ../RTL/cortexm0ds_logic.v(20231)
  // ../RTL/cortexm0ds_logic.v(18324)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4216|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6_reg  (
    .a({open_n33436,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykkiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 }),
    .mi({open_n33440,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 }),
    .f({_al_u4216_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykkiu6 }),
    .q({open_n33456,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 }));  // ../RTL/cortexm0ds_logic.v(18324)
  // ../RTL/cortexm0ds_logic.v(19715)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4217|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6_reg  (
    .b({_al_u4216_o,_al_u4219_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4217_o}),
    .f({_al_u4217_o,open_n33473}),
    .q({open_n33477,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 }));  // ../RTL/cortexm0ds_logic.v(19715)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4219|_al_u4218  (
    .a({open_n33478,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1600_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [4]}),
    .d({_al_u4218_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6]}),
    .f({_al_u4219_o,_al_u4218_o}));
  // ../RTL/cortexm0ds_logic.v(18192)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4222|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6_reg  (
    .a({open_n33499,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qgkiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 }),
    .mi({open_n33503,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .f({_al_u4222_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qgkiu6 }),
    .q({open_n33519,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 }));  // ../RTL/cortexm0ds_logic.v(18192)
  // ../RTL/cortexm0ds_logic.v(18975)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4223|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6_reg  (
    .b({_al_u4222_o,_al_u4225_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4223_o}),
    .f({_al_u4223_o,open_n33540}),
    .q({open_n33544,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 }));  // ../RTL/cortexm0ds_logic.v(18975)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4225|_al_u4224  (
    .a({open_n33545,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1592_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [2]}),
    .d({_al_u4224_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4]}),
    .f({_al_u4225_o,_al_u4224_o}));
  // ../RTL/cortexm0ds_logic.v(18191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4228|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6_reg  (
    .a({open_n33566,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0iiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 }),
    .mi({open_n33570,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .f({_al_u4228_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0iiu6 }),
    .q({open_n33586,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 }));  // ../RTL/cortexm0ds_logic.v(18191)
  // ../RTL/cortexm0ds_logic.v(18969)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4229|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6_reg  (
    .b({_al_u4228_o,_al_u4231_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4229_o}),
    .f({_al_u4229_o,open_n33607}),
    .q({open_n33611,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 }));  // ../RTL/cortexm0ds_logic.v(18969)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u422|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [1],\u_cmsdk_mcu/p1_out [1]}),
    .mi({open_n33615,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b1/B1_0 }),
    .q({open_n33630,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [1]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4231|_al_u4230  (
    .a({open_n33631,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({_al_u1573_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [3]}),
    .d({_al_u4230_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5]}),
    .f({_al_u4231_o,_al_u4230_o}));
  // ../RTL/cortexm0ds_logic.v(20186)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4234|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6_reg  (
    .a({open_n33656,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0niu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 }),
    .mi({open_n33667,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 }),
    .f({_al_u4234_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z0niu6 }),
    .q({open_n33672,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 }));  // ../RTL/cortexm0ds_logic.v(20186)
  // ../RTL/cortexm0ds_logic.v(17944)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(B*~(D*C*A))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(B*~(D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0100110011001100),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4235|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,open_n33673}),
    .b({_al_u4234_o,_al_u4237_o}),
    .c({_al_u1299_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 ,_al_u4235_o}),
    .f({_al_u4235_o,open_n33692}),
    .q({open_n33696,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 }));  // ../RTL/cortexm0ds_logic.v(17944)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4237|_al_u4236  (
    .a({open_n33697,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({_al_u3808_o,_al_u3797_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [8]}),
    .d({_al_u4236_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10]}),
    .f({_al_u4237_o,_al_u4236_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~C*~A*~(D*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000100000101),
    .MODE("LOGIC"))
    \_al_u4241|_al_u4240  (
    .a({_al_u4240_o,open_n33722}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Agyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .c({_al_u2296_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,_al_u1308_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 ,_al_u4240_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("~(A*~((D*B))*~(C)+A*(D*B)*~(C)+~(A)*(D*B)*C+A*(D*B)*C)"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0011010111110101),
    .MODE("LOGIC"))
    \_al_u4242|_al_u3386  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 ,open_n33743}),
    .b({_al_u1757_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kalpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .f({_al_u4242_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swyhu6 }));
  // ../RTL/cortexm0ds_logic.v(17576)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(D*~(C*~B))"),
    //.LUTG1("(D*~(C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000000),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1100111100000000),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4245|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6_reg  (
    .b({_al_u4244_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u2299_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .mi({open_n33769,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .f({_al_u4245_o,_al_u4244_o}),
    .q({open_n33785,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 }));  // ../RTL/cortexm0ds_logic.v(17576)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*C*~B))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1010101010001010),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u4246|_al_u3323  (
    .a({open_n33786,_al_u3322_o}),
    .b({open_n33787,_al_u3255_o}),
    .c({_al_u4244_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0zhu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 }),
    .f({_al_u4246_o,_al_u3323_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*~C*B))"),
    //.LUTF1("(D*~(C*~B*~A))"),
    //.LUTG0("(~A*~(D*~C*B))"),
    //.LUTG1("(D*~(C*~B*~A))"),
    .INIT_LUTF0(16'b0101000101010101),
    .INIT_LUTF1(16'b1110111100000000),
    .INIT_LUTG0(16'b0101000101010101),
    .INIT_LUTG1(16'b1110111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4248|_al_u4247  (
    .a({_al_u4245_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkzhu6 }),
    .b({_al_u4246_o,_al_u1251_o}),
    .c({_al_u4247_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .f({_al_u4248_o,_al_u4247_o}));
  // ../RTL/cortexm0ds_logic.v(17344)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(~D*~B)*~(C*~A))"),
    //.LUT1("(~C*B*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001110011),
    .INIT_LUT1(16'b0000110000000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4249|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6_reg  (
    .a({_al_u4239_o,_al_u4249_o}),
    .b({_al_u4243_o,_al_u1761_o}),
    .c({_al_u4248_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u4249_o,open_n33845}),
    .q({open_n33849,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }));  // ../RTL/cortexm0ds_logic.v(17344)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u424|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b10  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [10],\u_cmsdk_mcu/p1_out [10]}),
    .mi({open_n33853,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b10/B1_0 }),
    .q({open_n33868,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [10]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cortexm0ds_logic.v(20238)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(D*~A*~(C*B))"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(D*~A*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b0001010100000000),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b0001010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4251|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6_reg  (
    .a({_al_u3874_o,open_n33869}),
    .b({_al_u1774_o,open_n33870}),
    .c({_al_u1777_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ,_al_u4251_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4251_o,open_n33888}),
    .q({open_n33892,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 }));  // ../RTL/cortexm0ds_logic.v(20238)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u4254|_al_u1367  (
    .b({open_n33895,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }),
    .c({_al_u1367_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7cpw6_lutinv ,_al_u1367_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~C*~A*~(D*B))"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000100000101),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4256|_al_u4252  (
    .a({_al_u4252_o,_al_u4159_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7cpw6_lutinv ,_al_u679_o}),
    .c({_al_u4151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u4256_o,_al_u4252_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(D*C*~A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(D*C*~A))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000110011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4257|_al_u3124  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ,open_n33940}),
    .b({_al_u4256_o,open_n33941}),
    .c({_al_u3754_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u3124_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ,_al_u3124_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u4258|_al_u4255  (
    .a({open_n33966,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv ,_al_u1296_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,_al_u1344_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 ,_al_u2403_o}),
    .f({_al_u4258_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxaiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~D*~(C*B*A))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~D*~(C*B*A))"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0000000001111111),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0000000001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4260|_al_u3671  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv ,open_n33987}),
    .b({_al_u604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .c({_al_u1336_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u4259_o,_al_u1813_o}),
    .f({_al_u4260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwaiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~A*~(~D*~B)))"),
    //.LUTF1("(~D*~(C*~B*A))"),
    //.LUTG0("(C*~(~A*~(~D*~B)))"),
    //.LUTG1("(~D*~(C*~B*A))"),
    .INIT_LUTF0(16'b1010000010110000),
    .INIT_LUTF1(16'b0000000011011111),
    .INIT_LUTG0(16'b1010000010110000),
    .INIT_LUTG1(16'b0000000011011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4261|_al_u4345  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ,_al_u3085_o}),
    .b({_al_u4258_o,_al_u4344_o}),
    .c({_al_u4260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 }),
    .f({_al_u4261_o,_al_u4345_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("(C*~(B*D))"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"))
    \_al_u4263|_al_u4262  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .c({_al_u4262_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 }),
    .f({_al_u4263_o,_al_u4262_o}));
  // ../RTL/cortexm0ds_logic.v(17385)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*~B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4267|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6_reg  (
    .b({_al_u4266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y8lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u2299_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pyyhu6_lutinv }),
    .mi({open_n34070,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .f({_al_u4267_o,_al_u4266_o}),
    .q({open_n34075,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 }));  // ../RTL/cortexm0ds_logic.v(17385)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~A*~(~D*~C*B))"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~A*~(~D*~C*B))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0101010101010001),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4268|_al_u2305  (
    .a({_al_u2305_o,_al_u1757_o}),
    .b({_al_u2298_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jflpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yklpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2zhu6_lutinv ,_al_u2305_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~D*C*~B*A)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u4269|_al_u4243  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9zhu6 }),
    .b({_al_u4267_o,_al_u2295_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X2zhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A1zhu6_lutinv }),
    .d({_al_u3328_o,_al_u4242_o}),
    .f({_al_u4269_o,_al_u4243_o}));
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u426|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b11  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [11],\u_cmsdk_mcu/p1_out [11]}),
    .mi({open_n34123,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b11/B1_0 }),
    .q({open_n34138,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [11]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cortexm0ds_logic.v(17575)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*C*B))"),
    //.LUTF1("(D*~B*~(C*A))"),
    //.LUTG0("(A*~(~D*C*B))"),
    //.LUTG1("(D*~B*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000101010),
    .INIT_LUTF1(16'b0001001100000000),
    .INIT_LUTG0(16'b1010101000101010),
    .INIT_LUTG1(16'b0001001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4271|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .b({_al_u3390_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7zhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zslpw6 }),
    .mi({open_n34142,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .f({_al_u4271_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7zhu6 }),
    .q({open_n34158,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 }));  // ../RTL/cortexm0ds_logic.v(17575)
  // ../RTL/cortexm0ds_logic.v(17574)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*~C*A))"),
    //.LUT1("(D*~(~C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011000100),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4273|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6_reg  (
    .a({open_n34159,_al_u4239_o}),
    .b({_al_u4271_o,_al_u4273_o}),
    .c({_al_u4272_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u4269_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .mi({open_n34170,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }),
    .f({_al_u4273_o,_al_u4274_o}),
    .q({open_n34175,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 }));  // ../RTL/cortexm0ds_logic.v(17574)
  // ../RTL/cortexm0ds_logic.v(17350)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~B*~(~A*(D@C)))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~B*~(~A*(D@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0011001000100011),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0011001000100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4275|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6_reg  (
    .a({_al_u1761_o,open_n34176}),
    .b({_al_u1763_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1zhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bclpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 ,_al_u4274_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H1zhu6 ,open_n34194}),
    .q({open_n34198,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlpw6 }));  // ../RTL/cortexm0ds_logic.v(17350)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4277|_al_u7162  (
    .a({open_n34199,_al_u4289_o}),
    .b({open_n34200,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .d({_al_u4170_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [0]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr6ow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4278|_al_u4171  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 }),
    .d({_al_u4169_o,_al_u4170_o}),
    .f({_al_u4278_o,_al_u4171_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(D@B@A))"),
    //.LUTF1("(D*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    //.LUTG0("(C*(D@B@A))"),
    //.LUTG1("(D*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1001000001100000),
    .INIT_LUTF1(16'b1111110011000000),
    .INIT_LUTG0(16'b1001000001100000),
    .INIT_LUTG1(16'b1111110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4279|_al_u4421  (
    .a({open_n34249,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 }),
    .b({_al_u4278_o,_al_u4278_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ,_al_u3797_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0ghu6 ,_al_u4421_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*~(~A*~(D*B)))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1110000010100000),
    .MODE("LOGIC"))
    \_al_u4281|_al_u4280  (
    .a({_al_u4280_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv }),
    .b({_al_u2782_o,_al_u3690_o}),
    .c({_al_u696_o,_al_u604_o}),
    .d({_al_u3924_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 }),
    .f({_al_u4281_o,_al_u4280_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(B*~(D*~(~C*A)))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000100011001100),
    .MODE("LOGIC"))
    \_al_u4284|_al_u4283  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxaiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv }),
    .b({_al_u4282_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .c({_al_u4283_o,_al_u3924_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4284_o,_al_u4283_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4285|_al_u4299  (
    .c({\u_cmsdk_mcu/LOCKUPRESET ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u4284_o,_al_u4284_o}),
    .f({\u_cmsdk_mcu/n1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv }));
  // ../RTL/cmsdk_mcu_clkctrl.v(119)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4288|u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write ,\u_cmsdk_mcu/SYSRESETREQ }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/nxt_hrst ,\u_cmsdk_mcu/n1 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ,\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/nxt_hrst }),
    .q({open_n34362,\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg }));  // ../RTL/cmsdk_mcu_clkctrl.v(119)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u428|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b12  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [12],\u_cmsdk_mcu/p1_out [12]}),
    .mi({open_n34366,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b12/B1_0 }),
    .q({open_n34381,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [12]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u4290|_al_u7061  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ,_al_u4172_o}),
    .d({_al_u4172_o,_al_u4289_o}),
    .f({_al_u4290_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*~A))"),
    //.LUTF1("(A*~(B*~(~D*C)))"),
    //.LUTG0("(~(~D*B)*~(~C*~A))"),
    //.LUTG1("(A*~(B*~(~D*C)))"),
    .INIT_LUTF0(16'b1111101000110010),
    .INIT_LUTF1(16'b0010001010100010),
    .INIT_LUTG0(16'b1111101000110010),
    .INIT_LUTG1(16'b0010001010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4292|_al_u4291  (
    .a({_al_u4291_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u4292_o,_al_u4291_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4293|_al_u7192  (
    .a({_al_u4284_o,_al_u4289_o}),
    .b({_al_u4289_o,_al_u4290_o}),
    .c({_al_u4290_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] }),
    .d({_al_u4292_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [13]}),
    .f({_al_u4293_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eidow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~C*~B*~D)"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4296|_al_u4294  (
    .b({_al_u4294_o,_al_u1299_o}),
    .c({_al_u4295_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u4293_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nn8iu6 ,_al_u4294_o}));
  // ../RTL/cortexm0ds_logic.v(18561)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(~C*~(~B*~(~D*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b0000110000001110),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4297|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6_reg  (
    .a({_al_u4170_o,open_n34480}),
    .b({_al_u4278_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({_al_u4173_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u4297_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4297_o,open_n34494}),
    .q({open_n34498,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 }));  // ../RTL/cortexm0ds_logic.v(18561)
  // ../RTL/cortexm0ds_logic.v(17989)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(D*~B*~(~C*A))"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(D*~B*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b0011000100000000),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b0011000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4300|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6_reg  (
    .a({_al_u927_o,open_n34499}),
    .b({_al_u933_o,open_n34500}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ,_al_u4300_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4300_o,open_n34518}),
    .q({open_n34522,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 }));  // ../RTL/cortexm0ds_logic.v(17989)
  // ../RTL/cortexm0ds_logic.v(19727)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*(D@A)))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C*(D@A)))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111001110110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111001110110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4302|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 ,_al_u4170_o}),
    .b({_al_u3808_o,_al_u4302_o}),
    .c({_al_u1354_o,_al_u3797_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4302_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 }),
    .q({open_n34542,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 }));  // ../RTL/cortexm0ds_logic.v(19727)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4304|_al_u2399  (
    .a({open_n34543,_al_u678_o}),
    .b({_al_u678_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u4304_o,_al_u2399_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~A*~(C*B)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~(~A*~(C*B)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011101010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011101010),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4305|_al_u4306  (
    .a({open_n34568,_al_u4305_o}),
    .b({open_n34569,_al_u681_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sy2ju6 ,_al_u1342_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 }),
    .f({_al_u4305_o,_al_u4306_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*~C*B))"),
    //.LUTF1("(~B*A*~(D*C))"),
    //.LUTG0("(~A*~(D*~C*B))"),
    //.LUTG1("(~B*A*~(D*C))"),
    .INIT_LUTF0(16'b0101000101010101),
    .INIT_LUTF1(16'b0000001000100010),
    .INIT_LUTG0(16'b0101000101010101),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4309|_al_u4307  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8bow6 ,_al_u4306_o}),
    .b({_al_u4308_o,_al_u607_o}),
    .c({_al_u3201_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u4309_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8bow6 }));
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u430|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b13  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [13],\u_cmsdk_mcu/p1_out [13]}),
    .mi({open_n34621,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b13/B1_0 }),
    .q({open_n34636,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [13]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4310|_al_u3918  (
    .a({open_n34637,_al_u3666_o}),
    .b({open_n34638,_al_u3917_o}),
    .c({_al_u3917_o,_al_u909_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apaiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u4310_o,_al_u3918_o}));
  // ../RTL/cortexm0ds_logic.v(17753)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*~A))"),
    //.LUTF1("(D*~(B*~(C*~A)))"),
    //.LUTG0("(~(~D*C)*~(B*~A))"),
    //.LUTG1("(D*~(B*~(C*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1011101100001011),
    .INIT_LUTG1(16'b0111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4311|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6_reg  (
    .a({_al_u4304_o,_al_u4311_o}),
    .b({_al_u4309_o,_al_u4346_o}),
    .c({_al_u4310_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u696_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4311_o,open_n34680}),
    .q({open_n34684,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }));  // ../RTL/cortexm0ds_logic.v(17753)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4312|_al_u3607  (
    .c({_al_u2770_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({_al_u3211_o,_al_u3211_o}),
    .f({_al_u4312_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~D*C*A))"),
    //.LUT1("(A*~(D*C*B))"),
    .INIT_LUT0(16'b0011001100010011),
    .INIT_LUT1(16'b0010101010101010),
    .MODE("LOGIC"))
    \_al_u4315|_al_u4314  (
    .a({_al_u4314_o,_al_u4312_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 ,_al_u4313_o}),
    .c({_al_u2364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u4315_o,_al_u4314_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~D*C*~B*A)"),
    .INIT_LUT0(16'b1101001111011111),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u4317|_al_u4316  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vviiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 }),
    .b({_al_u4316_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({_al_u1269_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u4317_o,_al_u4316_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~C*~A*~(D*B))"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000100000101),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4319|_al_u4318  (
    .a({_al_u4312_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .b({_al_u3233_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 }),
    .c({_al_u4317_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({_al_u4318_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u4319_o,_al_u4318_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(D*C*A))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(D*C*A))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0001001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0001001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4321|_al_u4457  (
    .a({_al_u3211_o,open_n34773}),
    .b({_al_u4320_o,_al_u2367_o}),
    .c({_al_u2367_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,_al_u2364_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4bow6 ,_al_u4457_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(D*B)))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1101000001010000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u4323|_al_u4322  (
    .a({_al_u4315_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4bow6 }),
    .b({_al_u4319_o,_al_u3608_o}),
    .c({_al_u4322_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u4323_o,_al_u4322_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(A*~(~B*~(D*C)))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(A*~(~B*~(D*C)))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1010100010001000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1010100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4325|_al_u4324  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ,open_n34818}),
    .b({_al_u4324_o,_al_u2380_o}),
    .c({_al_u3902_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,_al_u2371_o}),
    .f({_al_u4325_o,_al_u4324_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(D*C)))"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b1010001000100010),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u4326|_al_u4327  (
    .a({open_n34843,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .b({_al_u1582_o,_al_u4326_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ,_al_u1342_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,_al_u2829_o}),
    .f({_al_u4326_o,_al_u4327_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~D*~(C*~B)))"),
    //.LUTF1("(~B*~(D*C*A))"),
    //.LUTG0("(~A*~(~D*~(C*~B)))"),
    //.LUTG1("(~B*~(D*C*A))"),
    .INIT_LUTF0(16'b0101010100010000),
    .INIT_LUTF1(16'b0001001100110011),
    .INIT_LUTG0(16'b0101010100010000),
    .INIT_LUTG1(16'b0001001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4329|_al_u4328  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .b({_al_u4328_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Frziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u4329_o,_al_u4328_o}));
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u432|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [14],\u_cmsdk_mcu/p1_out [14]}),
    .mi({open_n34891,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b14/B1_0 }),
    .q({open_n34906,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [14]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"))
    \_al_u4330|_al_u3223  (
    .a({_al_u3205_o,open_n34907}),
    .b({_al_u4327_o,open_n34908}),
    .c({_al_u4329_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({_al_u909_o,_al_u909_o}),
    .f({_al_u4330_o,_al_u3223_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(D*C))"),
    //.LUT1("(A*~(~D*C*B))"),
    .INIT_LUT0(16'b0000000100010001),
    .INIT_LUT1(16'b1010101000101010),
    .MODE("LOGIC"))
    \_al_u4333|_al_u4332  (
    .a({_al_u4332_o,_al_u3186_o}),
    .b({_al_u1346_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ,_al_u932_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv }),
    .f({_al_u4333_o,_al_u4332_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0101111100010011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0101111100010011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4334|_al_u4359  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L45iu6_lutinv }),
    .b({_al_u1269_o,_al_u682_o}),
    .c({_al_u1342_o,_al_u1342_o}),
    .d({_al_u1344_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u4334_o,_al_u4359_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4336|_al_u2645  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pu1ju6_lutinv ,open_n34975}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({_al_u4336_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(D*C*~B*A)"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4338|_al_u4337  (
    .a({_al_u4330_o,_al_u4334_o}),
    .b({_al_u4331_o,_al_u4336_o}),
    .c({_al_u4333_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv }),
    .d({_al_u4337_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u4338_o,_al_u4337_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"))
    \_al_u4340|_al_u3018  (
    .a({_al_u607_o,open_n35024}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,open_n35025}),
    .c({_al_u1346_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u4340_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf6ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~A*~(D*~B)))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(C*~(~A*~(D*~B)))"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1011000010100000),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1011000010100000),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4343|_al_u4342  (
    .a({open_n35046,_al_u930_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi7ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({_al_u4342_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4343_o,_al_u4342_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4344|_al_u4253  (
    .b({_al_u3624_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .d({_al_u4343_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ya1ju6_lutinv }),
    .f({_al_u4344_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpaow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~(~B*A)))"),
    //.LUT1("(~D*~C*B*A)"),
    .INIT_LUT0(16'b0010111100000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"))
    \_al_u4346|_al_u4341  (
    .a({_al_u4323_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 }),
    .b({_al_u4339_o,_al_u3109_o}),
    .c({_al_u4341_o,_al_u4340_o}),
    .d({_al_u4345_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4346_o,_al_u4341_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4348|_al_u7060  (
    .b({open_n35119,_al_u4289_o}),
    .c({_al_u1809_o,_al_u7059_o}),
    .d({_al_u4284_o,_al_u4284_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ,_al_u7060_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(~(D*~C)*~(~B*~A))"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(~(D*~C)*~(~B*~A))"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b1110000011101110),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b1110000011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4349|_al_u363  (
    .a({_al_u4278_o,open_n35144}),
    .b({_al_u4173_o,open_n35145}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgapw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4351|_al_u4352  (
    .b({open_n35172,_al_u678_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ,_al_u4351_o}),
    .f({_al_u4351_o,_al_u4352_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~A*~(~D*B)))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b1010000011100000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u4354|_al_u4353  (
    .a({_al_u1784_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 }),
    .b({_al_u4352_o,_al_u903_o}),
    .c({_al_u697_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({_al_u4353_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u4354_o,_al_u4353_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~D*~C*~B*A)"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"))
    \_al_u4356|_al_u4355  (
    .a({_al_u4354_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .b({_al_u4012_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .c({_al_u4283_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .d({_al_u4355_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4356_o,_al_u4355_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~B*~(~C*~D))"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0011001100110000),
    .MODE("LOGIC"))
    \_al_u4358|_al_u4167  (
    .b({_al_u1336_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u1643_o,_al_u1336_o}),
    .f({_al_u4358_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~C*~A*~(~D*~B))"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000010100000100),
    .MODE("LOGIC"))
    \_al_u4361|_al_u4360  (
    .a({_al_u3666_o,open_n35255}),
    .b({_al_u4359_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({_al_u4360_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv }),
    .f({_al_u4361_o,_al_u4360_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~A*~(D*B)))"),
    //.LUT1("(D*~(B*~(C*~A)))"),
    .INIT_LUT0(16'b0000111000001010),
    .INIT_LUT1(16'b0111001100000000),
    .MODE("LOGIC"))
    \_al_u4362|_al_u4331  (
    .a({_al_u4358_o,_al_u4016_o}),
    .b({_al_u4361_o,_al_u1806_o}),
    .c({_al_u1806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,_al_u3124_o}),
    .f({_al_u4362_o,_al_u4331_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(A*~(C*B)))"),
    //.LUTF1("(~(D*C)*~(B*A))"),
    //.LUTG0("(~D*~(A*~(C*B)))"),
    //.LUTG1("(~(D*C)*~(B*A))"),
    .INIT_LUTF0(16'b0000000011010101),
    .INIT_LUTF1(16'b0000011101110111),
    .INIT_LUTG0(16'b0000000011010101),
    .INIT_LUTG1(16'b0000011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4363|_al_u4364  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ,_al_u4363_o}),
    .b({_al_u607_o,_al_u4161_o}),
    .c({_al_u903_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 }),
    .d({_al_u2829_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u4363_o,_al_u4364_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*~A)"),
    //.LUT1("(~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000001000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"))
    \_al_u4365|_al_u4357  (
    .a({_al_u4356_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq3pw6_lutinv }),
    .b({_al_u4357_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I30ju6_lutinv }),
    .c({_al_u4362_o,_al_u1271_o}),
    .d({_al_u4364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 ,_al_u4357_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u4366|_al_u4980  (
    .a({open_n35340,_al_u4539_o}),
    .b({open_n35341,_al_u4912_o}),
    .c({_al_u4151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~D*~B*~A))"),
    //.LUT1("(C*~(B*~(D*~A)))"),
    .INIT_LUT0(16'b0000111100001110),
    .INIT_LUT1(16'b0111000000110000),
    .MODE("LOGIC"))
    \_al_u4367|_al_u4350  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dgapw6 ,_al_u4170_o}),
    .b({_al_u4350_o,_al_u4173_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 ,_al_u4168_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .f({_al_u4367_o,_al_u4350_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4368|_al_u4499  (
    .a({open_n35382,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphiu6_lutinv }),
    .b({open_n35383,_al_u4173_o}),
    .c({_al_u4367_o,_al_u4168_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ueapw6 }),
    .f({_al_u4368_o,_al_u4499_o}));
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u436|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2],open_n35404}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .mi({open_n35408,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [2],_al_u4587_o}),
    .q({open_n35423,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [2]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cortexm0ds_logic.v(18639)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4370|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ,_al_u4368_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3436 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 }),
    .q({open_n35443,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 }));  // ../RTL/cortexm0ds_logic.v(18639)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(B*~(D*~C*~A))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b1100100011001100),
    .MODE("LOGIC"))
    \_al_u4372|_al_u4371  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 ,open_n35444}),
    .b({_al_u4371_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y40ju6 }),
    .f({_al_u4372_o,_al_u4371_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u4374|_al_u4373  (
    .b({_al_u4373_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .d({_al_u3831_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({_al_u4374_o,_al_u4373_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4376|_al_u3416  (
    .b({open_n35489,_al_u3415_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .d({_al_u3997_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hm7ow6_lutinv }),
    .f({_al_u4376_o,_al_u3416_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~B*~(C*~A)))"),
    //.LUTF1("(C*~(~B*~(D*~A)))"),
    //.LUTG0("(D*~(~B*~(C*~A)))"),
    //.LUTG1("(C*~(~B*~(D*~A)))"),
    .INIT_LUTF0(16'b1101110000000000),
    .INIT_LUTF1(16'b1101000011000000),
    .INIT_LUTG0(16'b1101110000000000),
    .INIT_LUTG1(16'b1101000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4378|_al_u4377  (
    .a({_al_u4375_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 }),
    .b({_al_u4377_o,_al_u4376_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .f({_al_u4378_o,_al_u4377_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~C*~A*~(~D*B))"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000010100000001),
    .MODE("LOGIC"))
    \_al_u4381|_al_u4380  (
    .a({_al_u4379_o,_al_u604_o}),
    .b({_al_u2772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u4380_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u4381_o,_al_u4380_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4383|_al_u4382  (
    .b({_al_u682_o,_al_u3122_o}),
    .c({_al_u696_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .d({_al_u4382_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }),
    .f({_al_u4383_o,_al_u4382_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4384|_al_u2647  (
    .b({_al_u2392_o,open_n35586}),
    .c({_al_u2647_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u696_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u4384_o,_al_u2647_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~(C@B)))"),
    //.LUTF1("(~A*~(D*~C*B))"),
    //.LUTG0("(A*~(~D*~(C@B)))"),
    //.LUTG1("(~A*~(D*~C*B))"),
    .INIT_LUTF0(16'b1010101000101000),
    .INIT_LUTF1(16'b0101000101010101),
    .INIT_LUTG0(16'b1010101000101000),
    .INIT_LUTG1(16'b0101000101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4387|_al_u4386  (
    .a({_al_u4386_o,_al_u3246_o}),
    .b({_al_u908_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u4387_o,_al_u4386_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*A*~(D*B))"),
    //.LUT1("(D*C*B*~A)"),
    .INIT_LUT0(16'b0000001000001010),
    .INIT_LUT1(16'b0100000000000000),
    .MODE("LOGIC"))
    \_al_u4388|_al_u4385  (
    .a({_al_u4378_o,_al_u4383_o}),
    .b({_al_u4381_o,_al_u1812_o}),
    .c({_al_u4385_o,_al_u4384_o}),
    .d({_al_u4387_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u4388_o,_al_u4385_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"))
    \_al_u4389|_al_u4007  (
    .a({_al_u2369_o,open_n35655}),
    .b({_al_u4007_o,open_n35656}),
    .c({_al_u4373_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .f({_al_u4389_o,_al_u4007_o}));
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u438|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [3],\u_cmsdk_mcu/p1_out [3]}),
    .mi({open_n35680,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b3/B1_0 }),
    .q({open_n35695,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [3]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(B*~(A*~(D*~C)))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(B*~(A*~(D*~C)))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0100110001000100),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0100110001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4391|_al_u3090  (
    .a({_al_u4390_o,_al_u2386_o}),
    .b({_al_u2386_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxoiu6 }),
    .c({_al_u2380_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .f({_al_u4391_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjiow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u4394|_al_u4393  (
    .b({_al_u2364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyiiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({_al_u4393_o,_al_u2770_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia0ju6 ,_al_u4393_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u4395|_al_u4392  (
    .a({_al_u4392_o,open_n35742}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia0ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .c({_al_u2371_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wa0ju6 ,_al_u912_o}),
    .f({_al_u4395_o,_al_u4392_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*~(D*C*~B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*~(D*C*~B))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000101010101010),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4397|_al_u4335  (
    .a({_al_u4396_o,open_n35763}),
    .b({_al_u3109_o,open_n35764}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmjiu6_lutinv ,_al_u1266_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ,_al_u903_o}),
    .f({_al_u4397_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*C*~A))"),
    //.LUTF1("(A*~(D*C*~B))"),
    //.LUTG0("(~B*~(D*C*~A))"),
    //.LUTG1("(A*~(D*C*~B))"),
    .INIT_LUTF0(16'b0010001100110011),
    .INIT_LUTF1(16'b1000101010101010),
    .INIT_LUTG0(16'b0010001100110011),
    .INIT_LUTG1(16'b1000101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4398|_al_u3696  (
    .a({_al_u4397_o,_al_u3109_o}),
    .b({_al_u3109_o,_al_u696_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yljiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4398_o,_al_u3696_o}));
  // ../RTL/cortexm0ds_logic.v(17271)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*~A))"),
    //.LUTF1("(~C*~(B*~(D*~A)))"),
    //.LUTG0("(~(~D*C)*~(B*~A))"),
    //.LUTG1("(~C*~(B*~(D*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b1011101100001011),
    .INIT_LUTG1(16'b0000011100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4399|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6_reg  (
    .a({_al_u4372_o,_al_u4399_o}),
    .b({_al_u4398_o,_al_u4416_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u909_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4399_o,open_n35830}),
    .q({open_n35834,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }));  // ../RTL/cortexm0ds_logic.v(17271)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(B*~(~D*~C*~A))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1100110011001000),
    .MODE("LOGIC"))
    \_al_u4402|_al_u4401  (
    .a({_al_u4401_o,open_n35835}),
    .b({_al_u681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({_al_u3754_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u909_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqziu6 }),
    .f({_al_u4402_o,_al_u4401_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*~(~C*~B)))"),
    //.LUTF1("(C*A*~(D*B))"),
    //.LUTG0("(~A*~(D*~(~C*~B)))"),
    //.LUTG1("(C*A*~(D*B))"),
    .INIT_LUTF0(16'b0000000101010101),
    .INIT_LUTF1(16'b0010000010100000),
    .INIT_LUTG0(16'b0000000101010101),
    .INIT_LUTG1(16'b0010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4404|_al_u4403  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .b({_al_u4161_o,_al_u604_o}),
    .c({_al_u4403_o,_al_u679_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u4404_o,_al_u4403_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*~(C*~B)))"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b1010101000100000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u4405|_al_u4396  (
    .a({_al_u4402_o,_al_u4388_o}),
    .b({_al_u4404_o,_al_u4391_o}),
    .c({_al_u1643_o,_al_u4395_o}),
    .d({_al_u1635_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .f({_al_u4405_o,_al_u4396_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4408|_al_u4407  (
    .b({_al_u4407_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .d({_al_u3223_o,_al_u909_o}),
    .f({_al_u4408_o,_al_u4407_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(D*C))"),
    //.LUT1("(C*~(B*D))"),
    .INIT_LUT0(16'b0000000100010001),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"))
    \_al_u4409|_al_u4406  (
    .a({open_n35926,_al_u912_o}),
    .b({_al_u4408_o,_al_u2386_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .d({_al_u4406_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({_al_u4409_o,_al_u4406_o}));
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u440|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [4],\u_cmsdk_mcu/p1_out [4]}),
    .mi({open_n35950,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b4/B1_0 }),
    .q({open_n35965,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [4]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(B*~A*~(~D*C))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0100010000000100),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0100010000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4411|_al_u3574  (
    .a({_al_u4409_o,open_n35966}),
    .b({_al_u4410_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv }),
    .c({_al_u3574_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llaow6_lutinv }),
    .f({_al_u4411_o,_al_u3574_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(A)*~(D)+(C*B)*A*~(D)+~((C*B))*A*D+(C*B)*A*D)"),
    //.LUTF1("(C*B*~(~D*~A))"),
    //.LUTG0("~((C*B)*~(A)*~(D)+(C*B)*A*~(D)+~((C*B))*A*D+(C*B)*A*D)"),
    //.LUTG1("(C*B*~(~D*~A))"),
    .INIT_LUTF0(16'b0101010100111111),
    .INIT_LUTF1(16'b1100000010000000),
    .INIT_LUTG0(16'b0101010100111111),
    .INIT_LUTG1(16'b1100000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4412|_al_u4400  (
    .a({_al_u4400_o,_al_u3810_o}),
    .b({_al_u4405_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ia8iu6_lutinv }),
    .c({_al_u4411_o,_al_u909_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u4412_o,_al_u4400_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~(~B*~A))"),
    //.LUTF1("(A*~(D*~(~C*~B)))"),
    //.LUTG0("(D*C*~(~B*~A))"),
    //.LUTG1("(A*~(D*~(~C*~B)))"),
    .INIT_LUTF0(16'b1110000000000000),
    .INIT_LUTF1(16'b0000001010101010),
    .INIT_LUTG0(16'b1110000000000000),
    .INIT_LUTG1(16'b0000001010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4416|_al_u4415  (
    .a({_al_u4413_o,_al_u1812_o}),
    .b({_al_u4414_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({_al_u4415_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u4416_o,_al_u4415_o}));
  // ../RTL/cortexm0ds_logic.v(18435)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4419|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 ,open_n36041}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .clk(XTAL1_wire),
    .d({_al_u4368_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4419_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 }),
    .q({open_n36058,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jxgax6 }));  // ../RTL/cortexm0ds_logic.v(18435)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*B)*~(D*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0101000111110011),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u4423|_al_u4422  (
    .a({open_n36059,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3iiu6 }),
    .b({open_n36060,_al_u3808_o}),
    .c({_al_u4422_o,_al_u1581_o}),
    .d({_al_u4421_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3]}),
    .f({_al_u4423_o,_al_u4422_o}));
  // ../RTL/cortexm0ds_logic.v(18267)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4425|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6_reg  (
    .a({open_n36081,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4iiu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 }),
    .mi({open_n36092,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({_al_u4425_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4iiu6 }),
    .q({open_n36097,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 }));  // ../RTL/cortexm0ds_logic.v(18267)
  // ../RTL/cortexm0ds_logic.v(18968)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4426|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6_reg  (
    .b({_al_u4425_o,_al_u4426_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4423_o}),
    .f({_al_u4426_o,open_n36118}),
    .q({open_n36122,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 }));  // ../RTL/cortexm0ds_logic.v(18968)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u442|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [5],\u_cmsdk_mcu/p1_out [5]}),
    .mi({open_n36126,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b5/B1_0 }),
    .q({open_n36141,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [5]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cortexm0ds_logic.v(17818)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0011001100001111),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4436|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6_reg  (
    .a({open_n36142,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [4]}),
    .mi({open_n36146,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ,_al_u5830_o}),
    .q({open_n36162,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 }));  // ../RTL/cortexm0ds_logic.v(17818)
  // ../RTL/cortexm0ds_logic.v(18102)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4438|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ,_al_u5832_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .f({_al_u4438_o,open_n36179}),
    .q({open_n36183,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 }));  // ../RTL/cortexm0ds_logic.v(18102)
  // ../RTL/cmsdk_ahb_to_iop.v(96)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4445|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg1_b1  (
    .b({_al_u3797_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jc3pw6 }),
    .c({_al_u1888_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv }),
    .clk(XTAL1_wire),
    .d({_al_u4368_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jc3pw6 ,\u_cmsdk_mcu/HSIZE [1]}),
    .q({open_n36206,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [1]}));  // ../RTL/cmsdk_ahb_to_iop.v(96)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(B*~(~D*~C)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~A*~(B*~(~D*~C)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0001000100010101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001000100010101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4448|_al_u526  (
    .a({open_n36207,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 }),
    .b({open_n36208,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gnqpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ,_al_u526_o}));
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u444|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6],open_n36233}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6],open_n36234}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n246 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [6],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [6],open_n36251}),
    .q({open_n36255,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [6]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cortexm0ds_logic.v(18101)
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    //.LUT1("(~D*C*B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111111),
    .INIT_LUT1(16'b0000000001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4450|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,open_n36256}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 ,open_n36257}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ,open_n36258}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 }),
    .mi({open_n36269,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({_al_u4450_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 }),
    .q({open_n36274,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 }));  // ../RTL/cortexm0ds_logic.v(18101)
  // ../RTL/cortexm0ds_logic.v(18219)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*B))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4451|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zrhiu6_lutinv ,_al_u4451_o}),
    .b({_al_u1777_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 }),
    .c({_al_u3925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u4450_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 }),
    .mi({open_n36285,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .f({_al_u4451_o,_al_u4452_o}),
    .q({open_n36290,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 }));  // ../RTL/cortexm0ds_logic.v(18219)
  // ../RTL/cortexm0ds_logic.v(18176)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4455|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6_reg  (
    .a({open_n36291,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfliu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 }),
    .mi({open_n36302,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .f({_al_u4455_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfliu6 }),
    .q({open_n36307,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 }));  // ../RTL/cortexm0ds_logic.v(18176)
  // ../RTL/cortexm0ds_logic.v(19729)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D*C*A))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011001100110011),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4456|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6_reg  (
    .a({open_n36308,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 }),
    .b({_al_u4455_o,_al_u4456_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ql8iu6 ,_al_u4457_o}),
    .f({_al_u4456_o,open_n36323}),
    .q({open_n36327,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 }));  // ../RTL/cortexm0ds_logic.v(19729)
  // ../RTL/cortexm0ds_logic.v(19557)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4459|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2phu6 ,open_n36328}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxdpw6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bggiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ,_al_u3339_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4459_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxdpw6 }),
    .q({open_n36349,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 }));  // ../RTL/cortexm0ds_logic.v(19557)
  // ../RTL/cortexm0ds_logic.v(19389)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4460|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W1phu6 ,open_n36350}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0phu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ,_al_u3468_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ,_al_u3467_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4460_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0phu6 }),
    .q({open_n36371,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 }));  // ../RTL/cortexm0ds_logic.v(19389)
  // ../RTL/cortexm0ds_logic.v(19449)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4461|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szohu6 ,open_n36372}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwdpw6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ,_al_u3489_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ,_al_u3488_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4461_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Szohu6 }),
    .q({open_n36393,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 }));  // ../RTL/cortexm0ds_logic.v(19449)
  // ../RTL/cortexm0ds_logic.v(19377)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4462|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B1phu6 ,open_n36394}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdpw6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ,_al_u3463_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ,_al_u3462_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4462_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B1phu6 }),
    .q({open_n36411,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 }));  // ../RTL/cortexm0ds_logic.v(19377)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u4463|_al_u6520  (
    .a({_al_u4459_o,open_n36412}),
    .b({_al_u4460_o,open_n36413}),
    .c({_al_u4461_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 }),
    .d({_al_u4462_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 }),
    .f({_al_u4463_o,_al_u6520_o}));
  // ../RTL/cortexm0ds_logic.v(20031)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4464|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F3phu6 ,open_n36434}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzohu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbdiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ,_al_u3483_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4464_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zzohu6 }),
    .q({open_n36451,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 }));  // ../RTL/cortexm0ds_logic.v(20031)
  // ../RTL/cortexm0ds_logic.v(19425)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4465|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0phu6 ,open_n36452}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0phu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ,_al_u3479_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ,_al_u3478_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4465_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0phu6 }),
    .q({open_n36469,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 }));  // ../RTL/cortexm0ds_logic.v(19425)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4466|_al_u6526  (
    .b({_al_u4464_o,open_n36472}),
    .c({_al_u4465_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 }),
    .d({_al_u4463_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 }),
    .f({_al_u4466_o,_al_u6526_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4467|_al_u6630  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 ,open_n36499}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 }),
    .d({_al_u4466_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 }),
    .f({_al_u4467_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17199)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~C*~B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111110001010100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4468|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jyohu6 ,open_n36524}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qh5iu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ,_al_u3520_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ,_al_u3519_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4468_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jyohu6 }),
    .q({open_n36541,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 }));  // ../RTL/cortexm0ds_logic.v(17199)
  // ../RTL/cortexm0ds_logic.v(19533)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4469|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4phu6 ,open_n36542}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4phu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ,_al_u3281_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ,_al_u3279_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux5iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4phu6 }),
    .q({open_n36559,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 }));  // ../RTL/cortexm0ds_logic.v(19533)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u446|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [7],\u_cmsdk_mcu/p1_out [7]}),
    .mi({open_n36563,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b7/B1_0 }),
    .q({open_n36578,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [7]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cortexm0ds_logic.v(19545)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(B*~(~C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4470|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux5iu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ,_al_u3372_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3phu6 ,_al_u3371_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4470_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3phu6 }),
    .q({open_n36597,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 }));  // ../RTL/cortexm0ds_logic.v(19545)
  // ../RTL/cortexm0ds_logic.v(19521)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(C*A*~(~D*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(C*A*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1010000000100000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1010000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4471|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6_reg  (
    .a({_al_u4468_o,open_n36598}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cyohu6 ,_al_u1777_o}),
    .c({_al_u4470_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Webiu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ,_al_u3524_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4471_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cyohu6 }),
    .q({open_n36619,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 }));  // ../RTL/cortexm0ds_logic.v(19521)
  // ../RTL/cortexm0ds_logic.v(19830)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4472|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3phu6 ,open_n36620}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1phu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9fiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ,_al_u3361_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4472_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3phu6 }),
    .q({open_n36637,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 }));  // ../RTL/cortexm0ds_logic.v(19830)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~C*B*~D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4473|_al_u5068  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv ,_al_u5067_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 }),
    .d({_al_u2733_o,_al_u5066_o}),
    .f({_al_u4473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 }));
  // ../RTL/cortexm0ds_logic.v(19281)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~B*~(~C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4474|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6_reg  (
    .b({_al_u4473_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ,_al_u3335_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5phu6 ,_al_u3334_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4474_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5phu6 }),
    .q({open_n36686,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 }));  // ../RTL/cortexm0ds_logic.v(19281)
  // ../RTL/cortexm0ds_logic.v(19365)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(~C*B)*~(~D*~A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(~C*B)*~(~D*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111001110100010),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111001110100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4475|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 ,open_n36687}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P1phu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ,_al_u3535_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4475_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P1phu6 }),
    .q({open_n36708,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 }));  // ../RTL/cortexm0ds_logic.v(19365)
  // ../RTL/cortexm0ds_logic.v(19401)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(B*A*~(~D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1000100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4476|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6_reg  (
    .a({_al_u4474_o,open_n36709}),
    .b({_al_u4475_o,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5phu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ,_al_u3457_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5phu6 }),
    .q({open_n36726,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 }));  // ../RTL/cortexm0ds_logic.v(19401)
  // ../RTL/cortexm0ds_logic.v(20144)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4477|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4phu6 ,open_n36727}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V4phu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ,_al_u3271_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ,_al_u3268_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O16iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4phu6 }),
    .q({open_n36744,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 }));  // ../RTL/cortexm0ds_logic.v(20144)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4478|_al_u6516  (
    .b({_al_u4476_o,open_n36747}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O16iu6 ,_al_u6510_o}),
    .d({_al_u4472_o,_al_u6509_o}),
    .f({_al_u4478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L3sow6_lutinv }));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000001110111),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b0010000001110111),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4479|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K2phu6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2phu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 }),
    .mi({open_n36775,\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vu5iu6 ,_al_u3352_o}),
    .q({open_n36790,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [14]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000001110111),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4480|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b9  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2phu6 ,\u_cmsdk_mcu/HWDATA [9]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwdpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 }),
    .mi({open_n36801,\u_cmsdk_mcu/HWDATA [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4480_o,_al_u3286_o}),
    .q({open_n36805,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [9]}));  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4481|_al_u5124  (
    .a({_al_u4471_o,open_n36806}),
    .b({_al_u4478_o,open_n36807}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vu5iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgeow6 }),
    .d({_al_u4480_o,_al_u5031_o}),
    .f({_al_u4481_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 }));
  // ../RTL/cortexm0ds_logic.v(19485)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4482|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzohu6 ,open_n36832}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezohu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfiu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ,_al_u3509_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zi5iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ezohu6 }),
    .q({open_n36853,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 }));  // ../RTL/cortexm0ds_logic.v(19485)
  // ../RTL/cortexm0ds_logic.v(19509)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4483|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xyohu6 ,open_n36854}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyohu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ,_al_u3530_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ,_al_u3529_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4483_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyohu6 }),
    .q({open_n36871,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 }));  // ../RTL/cortexm0ds_logic.v(19509)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4484|_al_u6449  (
    .a({_al_u4467_o,open_n36872}),
    .b({_al_u4481_o,open_n36873}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zi5iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 }),
    .d({_al_u4483_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 }),
    .f({_al_u4484_o,_al_u6449_o}));
  // ../RTL/cortexm0ds_logic.v(18993)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(C*~(A*~(~D*B)))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(C*~(A*~(~D*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0101000011010000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0101000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4485|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6_reg  (
    .a({_al_u4484_o,open_n36898}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npghu6 ,_al_u1777_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 ,_al_u1791_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ,_al_u3875_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4485_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npghu6 }),
    .q({open_n36919,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 }));  // ../RTL/cortexm0ds_logic.v(18993)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~D*~B*~(C*A))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~D*~B*~(C*A))"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0000000000010011),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0000000000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4487|_al_u4486  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwcpw6_lutinv ,open_n36920}),
    .b({_al_u3925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({_al_u4486_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv }),
    .f({_al_u4487_o,_al_u4486_o}));
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u448|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b8  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [8],\u_cmsdk_mcu/p1_out [8]}),
    .mi({open_n36948,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b8/B1_0 }),
    .q({open_n36963,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [8]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cortexm0ds_logic.v(18429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~B*~(~C*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0011001100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4490|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u4419_o,_al_u4419_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4490_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .q({open_n36981,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }));  // ../RTL/cortexm0ds_logic.v(18429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4491|_al_u4537  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ,open_n36984}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .d({_al_u4490_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 ,_al_u4537_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4493|_al_u4435  (
    .b({_al_u4492_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 }));
  // ../RTL/cortexm0ds_logic.v(18378)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4494|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bqzhu6_lutinv ,open_n37037}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 }),
    .mi({open_n37048,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n265 }),
    .q({open_n37052,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 }));  // ../RTL/cortexm0ds_logic.v(18378)
  // ../RTL/cortexm0ds_logic.v(18412)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(D*C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4495|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ,open_n37053}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 ,_al_u4197_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .mi({open_n37064,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .f({_al_u4495_o,_al_u4545_o}),
    .q({open_n37069,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 }));  // ../RTL/cortexm0ds_logic.v(18412)
  // ../RTL/cortexm0ds_logic.v(18724)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~B*~(~D*~(C*A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0011001100100000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4498|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6_reg  (
    .a({_al_u4171_o,open_n37070}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,open_n37071}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 ,_al_u4173_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,_al_u4171_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphiu6_lutinv ,open_n37084}),
    .q({open_n37088,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 }));  // ../RTL/cortexm0ds_logic.v(18724)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4500|_al_u4502  (
    .c({_al_u4499_o,_al_u4501_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aphiu6 ,_al_u4500_o}),
    .f({_al_u4500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4501|_al_u4048  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED ,open_n37113}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jcpow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED }),
    .f({_al_u4501_o,_al_u4048_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4504|_al_u4503  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ,_al_u1299_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17793)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(~D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111011111110111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4505|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu8iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,_al_u4509_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ,_al_u4530_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu8iu6 ,open_n37179}),
    .q({open_n37183,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }));  // ../RTL/cortexm0ds_logic.v(17793)
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*~(~D*B))"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1010000000100000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u4506|_al_u4510  (
    .a({open_n37184,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(A*~(~D*B)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000010100001101),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4508|_al_u4507  (
    .a({open_n37205,_al_u4170_o}),
    .b({open_n37206,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ekhiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8jax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vihiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ekhiu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(20213)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*~D))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~C*~(B*~D))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000011111100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4509|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ,open_n37227}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6 ,_al_u1286_o}),
    .f({_al_u4509_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw8iu6 }),
    .q({open_n37248,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Swjbx6 }));  // ../RTL/cortexm0ds_logic.v(20213)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b0010010110100001),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b0010010110100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u450|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b9  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [9],\u_cmsdk_mcu/p1_out [9]}),
    .mi({open_n37252,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b9/B1_0 }),
    .q({open_n37267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [9]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4512|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b14  (
    .a({_al_u1986_o,open_n37268}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n37269}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n181 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n217 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [14],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4512_o,open_n37286}),
    .q({open_n37290,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [14]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4513|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n37291}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n37292}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n226 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n262 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [14],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4513_o,open_n37309}),
    .q({open_n37313,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [14]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(~D*C))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~B*~A*~(~D*C))"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0001000100000001),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0001000100000001),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4514|_al_u4577  (
    .a({open_n37314,_al_u4574_o}),
    .b({_al_u1982_o,_al_u4575_o}),
    .c({_al_u4513_o,_al_u1982_o}),
    .d({_al_u4512_o,_al_u4576_o}),
    .f({_al_u4514_o,_al_u4577_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4516|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n37339}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n37340}),
    .c({\u_cmsdk_mcu/p0_outen [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n82 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [14],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4516_o,open_n37353}),
    .q({open_n37357,\u_cmsdk_mcu/p0_outen [14]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b0011000100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4517|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b14  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [14]}),
    .b({_al_u4516_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [14],\u_cmsdk_mcu/p0_out [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4517_o,open_n37370}),
    .q({open_n37374,\u_cmsdk_mcu/p0_out [14]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4518|_al_u4825  (
    .a({_al_u4511_o,_al_u4511_o}),
    .b({_al_u4514_o,_al_u4822_o}),
    .c({_al_u4517_o,_al_u4824_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [8]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4519|_al_u4828  (
    .a({_al_u1986_o,_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [8]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [8]}),
    .f({_al_u4519_o,_al_u4828_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b1000101111001111),
    .MODE("LOGIC"))
    \_al_u4520|_al_u4806  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [12]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[12] }),
    .f({_al_u4520_o,_al_u4806_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4521|_al_u4731  (
    .b({_al_u1982_o,_al_u1982_o}),
    .c({_al_u4520_o,_al_u4730_o}),
    .d({_al_u4519_o,_al_u4729_o}),
    .f({_al_u4521_o,_al_u4731_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4523|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n37469}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n37470}),
    .c({\u_cmsdk_mcu/p1_outen [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n46 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n82 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [14],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4523_o,open_n37483}),
    .q({open_n37487,\u_cmsdk_mcu/p1_outen [14]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*~(~B*~(~C*A)))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*~(~B*~(~C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011001110),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4524|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b14/B1_0 ,open_n37488}),
    .b({_al_u4523_o,open_n37489}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/p1_outen [14]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/p1_out [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4524_o,open_n37507}),
    .q({open_n37511,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [14]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~D*~(A*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000000001011101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4526|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4521_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4524_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]}),
    .clk(XTAL1_wire),
    .d({_al_u4525_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]}),
    .mi({open_n37523,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4526_o,_al_u4525_o}),
    .q({open_n37527,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [14]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4528|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b14  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n37528}),
    .b({_al_u4527_o,open_n37529}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [14]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4528_o,open_n37546}),
    .q({open_n37550,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [14]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u452|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b3  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [3],open_n37553}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u452_o,open_n37566}),
    .q({open_n37570,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [3]}));  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(D*~A))"),
    //.LUT1("(~C*~(B*~D))"),
    .INIT_LUT0(16'b1000000011000000),
    .INIT_LUT1(16'b0000111100000011),
    .MODE("LOGIC"))
    \_al_u4530|_al_u6725  (
    .a({open_n37571,_al_u4529_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ,_al_u6722_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ,_al_u6724_o}),
    .d({_al_u4529_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u4530_o,_al_u6725_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u4533|_al_u6744  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ,_al_u4533_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv ,_al_u6743_o}),
    .f({_al_u4533_o,_al_u6744_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~D))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0011001100000011),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u4534|_al_u4532  (
    .b({_al_u4532_o,_al_u4501_o}),
    .c({_al_u4533_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ,_al_u4500_o}),
    .f({_al_u4534_o,_al_u4532_o}));
  // ../RTL/cortexm0ds_logic.v(18645)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4535|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 ,open_n37638}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,open_n37639}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vobiu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4535_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .q({open_n37659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tajax6 }));  // ../RTL/cortexm0ds_logic.v(18645)
  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u453|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg5_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [0],open_n37662}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .clk(XTAL1_wire),
    .d({_al_u452_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u453_o,open_n37679}),
    .q({open_n37683,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [1]}));  // ../RTL/cmsdk_apb_uart.v(405)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4540|_al_u4539  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iiliu6 ,_al_u1888_o}),
    .d({_al_u4539_o,_al_u4368_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ,_al_u4539_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4542|_al_u2272  (
    .a({open_n37712,_al_u1888_o}),
    .b({_al_u3797_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qk9pw6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8lax6 }),
    .d({_al_u4539_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .f({_al_u4542_o,_al_u2272_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4544|_al_u4496  (
    .b({_al_u3887_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 ,_al_u4495_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u4544_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4548|_al_u4547  (
    .a({_al_u4544_o,open_n37763}),
    .b({_al_u4545_o,_al_u4101_o}),
    .c({_al_u4546_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u4548_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv }));
  // ../RTL/cortexm0ds_logic.v(18044)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4549|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6_reg  (
    .a({open_n37788,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [10]}),
    .mi({open_n37792,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .f({_al_u4549_o,_al_u5818_o}),
    .q({open_n37808,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 }));  // ../RTL/cortexm0ds_logic.v(18044)
  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~B*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111111111111100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111111111111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u454|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b6  (
    .b({_al_u453_o,open_n37811}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [6],_al_u2488_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n53 ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n37815,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n246 }),
    .q({open_n37830,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [6]}));  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    //.LUT1("(~A*~(~B*~(D*C)))"),
    .INIT_LUT0(16'b0010000010101000),
    .INIT_LUT1(16'b0101010001000100),
    .MODE("LOGIC"))
    \_al_u4552|_al_u4916  (
    .a({_al_u4550_o,_al_u4552_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .c({_al_u4551_o,_al_u4086_o}),
    .d({_al_u4091_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 }),
    .f({_al_u4552_o,_al_u4916_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4556|_al_u4555  (
    .c({_al_u4533_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz4iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 }));
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4557|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b1  (
    .a({_al_u1986_o,open_n37875}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n37876}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n191 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4557_o,open_n37889}),
    .q({open_n37893,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [1]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000101111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4558|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n37894}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n37895}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n236 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4558_o,open_n37908}),
    .q({open_n37912,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [1]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4559|_al_u4703  (
    .b({_al_u1982_o,_al_u1982_o}),
    .c({_al_u4558_o,_al_u4702_o}),
    .d({_al_u4557_o,_al_u4701_o}),
    .f({_al_u4559_o,_al_u4703_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4560|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n37935}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n37936}),
    .c({\u_cmsdk_mcu/p0_outen [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n56 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4560_o,open_n37953}),
    .q({open_n37957,\u_cmsdk_mcu/p0_outen [1]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4561|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b1  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [1]}),
    .b({_al_u4560_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4:3]),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [1],\u_cmsdk_mcu/p0_out [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4561_o,open_n37974}),
    .q({open_n37978,\u_cmsdk_mcu/p0_out [1]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u4562|_al_u4785  (
    .a({_al_u4511_o,_al_u4511_o}),
    .b({_al_u4559_o,_al_u4782_o}),
    .c({_al_u4561_o,_al_u4784_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4562_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [11]}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110101011000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4564|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({_al_u4563_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4564_o,open_n38011}),
    .q({open_n38015,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [1]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4568|_al_u4567  (
    .a({_al_u4562_o,_al_u1988_o}),
    .b({_al_u4564_o,_al_u1986_o}),
    .c({_al_u4567_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],_al_u4566_o}),
    .f({_al_u4568_o,_al_u4567_o}));
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u456|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b13  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2],_al_u4136_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u456_o,\u_cmsdk_mcu/HADDR [15]}),
    .q({open_n38057,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [15]}));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4570|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b5  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .clk(XTAL1_wire),
    .d({_al_u4569_o,_al_u496_o}),
    .mi({open_n38070,\u_cmsdk_mcu/HADDR [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ,_al_u497_o}),
    .q({open_n38074,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [7]}));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4571|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg2_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ,open_n38075}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [1],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .f({_al_u4571_o,open_n38088}),
    .q({open_n38092,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [1]}));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4573|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38093}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/p1_outen [1]}),
    .c({\u_cmsdk_mcu/p1_outen [1],\u_cmsdk_mcu/p1_altfunc [1]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [1],\u_cmsdk_mcu/p1_out [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4573_o,open_n38107}),
    .q({open_n38111,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [1]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~B*~(~C*A)))"),
    //.LUTF1("(~D*~(~B*~(~C*A)))"),
    //.LUTG0("(~D*~(~B*~(~C*A)))"),
    //.LUTG1("(~D*~(~B*~(~C*A)))"),
    .INIT_LUTF0(16'b0000000011001110),
    .INIT_LUTF1(16'b0000000011001110),
    .INIT_LUTG0(16'b0000000011001110),
    .INIT_LUTG1(16'b0000000011001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4574|_al_u4872  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b1/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b13/B1_0 }),
    .b({_al_u4573_o,_al_u4871_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4574_o,_al_u4872_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"))
    \_al_u4575|_al_u4788  (
    .a({_al_u1986_o,_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [11]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [11]}),
    .f({_al_u4575_o,_al_u4788_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4576|_al_u4754  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [9]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[9] }),
    .f({_al_u4576_o,_al_u4754_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*B))"),
    //.LUT1("(D*~(C*~(~B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b0010111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4579|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,_al_u4567_o}),
    .b({_al_u4577_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .c({_al_u4578_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]}),
    .mi({open_n38191,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [1],_al_u4578_o}),
    .q({open_n38195,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [1]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000001000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u457|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b10  (
    .a({_al_u456_o,open_n38196}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [12],_al_u4035_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 ,\u_cmsdk_mcu/HADDR [12]}),
    .q({open_n38212,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [12]}));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4580|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable ,\u_cmsdk_mcu/HWRITE }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4580_o,open_n38233}),
    .q({open_n38237,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_read_enable }));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  // ../RTL/cortexm0ds_logic.v(17417)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4582|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,_al_u4582_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,_al_u4584_o}),
    .c({_al_u4581_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1833_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4582_o,open_n38251}),
    .q({open_n38255,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }));  // ../RTL/cortexm0ds_logic.v(17417)
  // ../RTL/cortexm0ds_logic.v(18223)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010111000111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4584|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6_reg  (
    .a({open_n38256,_al_u4500_o}),
    .b({_al_u4583_o,_al_u4501_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7mpw6 }),
    .mi({open_n38267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .f({_al_u4584_o,_al_u4583_o}),
    .q({open_n38272,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 }));  // ../RTL/cortexm0ds_logic.v(18223)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*C*~D+~A*~B*C*D+~A*B*C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4586|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b2_rom0  (
    .a({open_n38273,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4586_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b1000101111001111),
    .MODE("LOGIC"))
    \_al_u4588|_al_u4680  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [5]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[5] }),
    .f({_al_u4588_o,_al_u4680_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4591|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38314}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n38315}),
    .c({\u_cmsdk_mcu/p1_outen [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4591_o,open_n38328}),
    .q({open_n38332,\u_cmsdk_mcu/p1_outen [2]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~B*~(~C*A)))"),
    //.LUTF1("(~D*~(~B*~(~C*A)))"),
    //.LUTG0("(~D*~(~B*~(~C*A)))"),
    //.LUTG1("(~D*~(~B*~(~C*A)))"),
    .INIT_LUTF0(16'b0000000011001110),
    .INIT_LUTF1(16'b0000000011001110),
    .INIT_LUTG0(16'b0000000011001110),
    .INIT_LUTG1(16'b0000000011001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4592|_al_u4858  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b2/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b0/B1_0 }),
    .b({_al_u4591_o,_al_u4857_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4592_o,_al_u4858_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4593|_al_u4768  (
    .a({_al_u1986_o,_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [10]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [10]}),
    .f({_al_u4593_o,_al_u4768_o}));
  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(D*~(C*B)))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(~A*~(D*~(C*B)))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111110101010),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1011111110101010),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4595|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg2_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ,\u_cmsdk_mcu/n1 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ,\u_cmsdk_mcu/HWDATA [2]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .f({_al_u4595_o,open_n38397}),
    .q({open_n38401,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [2]}));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4596|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b2  (
    .a({_al_u1986_o,open_n38402}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38403}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n193 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4596_o,open_n38420}),
    .q({open_n38424,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [2]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000101111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4597|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n38425}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38426}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n238 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4597_o,open_n38439}),
    .q({open_n38443,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [2]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4598|_al_u4684  (
    .b({_al_u1982_o,_al_u1982_o}),
    .c({_al_u4597_o,_al_u4683_o}),
    .d({_al_u4596_o,_al_u4682_o}),
    .f({_al_u4598_o,_al_u4684_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4599|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38466}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n38467}),
    .c({\u_cmsdk_mcu/p0_outen [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [2],\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4599_o,open_n38480}),
    .q({open_n38484,\u_cmsdk_mcu/p0_outen [2]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_ahb_to_apb.v(253)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(D*A*(C@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0010100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u459|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg2_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],open_n38485}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n43 ,open_n38499}),
    .q({open_n38503,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]}));  // ../RTL/cmsdk_ahb_to_apb.v(253)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b0011000100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4600|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b2  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [2]}),
    .b({_al_u4599_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [2],\u_cmsdk_mcu/p0_out [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4600_o,open_n38516}),
    .q({open_n38520,\u_cmsdk_mcu/p0_out [2]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4602|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b8  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [8],_al_u4111_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u4602_o,\u_cmsdk_mcu/HADDR [10]}),
    .q({open_n38539,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [8]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4603|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b6  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [5],_al_u4106_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({_al_u4602_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u4603_o,\u_cmsdk_mcu/HADDR [8]}),
    .q({open_n38562,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [6]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4604|_al_u4667  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]}),
    .d({_al_u4603_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [4]}),
    .f({_al_u4604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [5]}));
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4605|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8],open_n38591}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2],_al_u4219_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u4605_o,\u_cmsdk_mcu/HADDR [5]}),
    .q({open_n38612,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*(D@C))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*A*(D@C))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000100010000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4606|_al_u4632  (
    .a({open_n38613,_al_u4604_o}),
    .b({open_n38614,_al_u4631_o}),
    .c({_al_u4605_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1]}),
    .d({_al_u4604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [3]}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*C)*~(B*A))"),
    //.LUTG0("~(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110101011000000),
    .INIT_LUTF1(16'b0000011101110111),
    .INIT_LUTG0(16'b1110101011000000),
    .INIT_LUTG1(16'b0000011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4607|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b2  (
    .a({\u_cmsdk_mcu/sram_hrdata [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4607_o,open_n38655}),
    .q({open_n38659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [2]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4608|_al_u4635  (
    .a({open_n38660,_al_u4633_o}),
    .b({\u_cmsdk_mcu/flash_hrdata [2],_al_u4634_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/sram_hrdata [3]}),
    .d({_al_u4607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}),
    .f({_al_u4608_o,_al_u4635_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4609|_al_u4511  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [2],open_n38681}),
    .b({_al_u4586_o,open_n38682}),
    .c({_al_u4608_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o }),
    .f({_al_u4609_o,_al_u4511_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(C*~B*~(D*~A))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(C*~B*~(D*~A))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0010000000110000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0010000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4610|_al_u4601  (
    .a({_al_u4595_o,_al_u4511_o}),
    .b({_al_u4601_o,_al_u4598_o}),
    .c({_al_u4609_o,_al_u4600_o}),
    .d({_al_u4580_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4610_o,_al_u4601_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4611|_al_u4594  (
    .a({open_n38731,_al_u4589_o}),
    .b({_al_u4610_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],_al_u4592_o}),
    .d({_al_u4594_o,_al_u4593_o}),
    .f({_al_u4611_o,_al_u4594_o}));
  // ../RTL/cortexm0ds_logic.v(17442)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4612|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,_al_u4612_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uehiu6 }),
    .c({_al_u4611_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1836_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4612_o,open_n38769}),
    .q({open_n38773,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }));  // ../RTL/cortexm0ds_logic.v(17442)
  // ../RTL/cortexm0ds_logic.v(18193)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010111000111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4614|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6_reg  (
    .a({open_n38774,_al_u4500_o}),
    .b({_al_u4613_o,_al_u4501_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 }),
    .mi({open_n38785,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uehiu6 ,_al_u4613_o}),
    .q({open_n38790,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 }));  // ../RTL/cortexm0ds_logic.v(18193)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4616|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b3  (
    .a({_al_u1986_o,open_n38791}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38792}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n195 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4616_o,open_n38805}),
    .q({open_n38809,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [3]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4617|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n38810}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38811}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n240 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4617_o,open_n38828}),
    .q({open_n38832,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [3]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4618|_al_u4644  (
    .b({_al_u1982_o,_al_u1982_o}),
    .c({_al_u4617_o,_al_u4643_o}),
    .d({_al_u4616_o,_al_u4642_o}),
    .f({_al_u4618_o,_al_u4644_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4619|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38859}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n38860}),
    .c({\u_cmsdk_mcu/p0_outen [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n60 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4619_o,open_n38877}),
    .q({open_n38881,\u_cmsdk_mcu/p0_outen [3]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4620|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b3  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [3]}),
    .b({_al_u4619_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [3],\u_cmsdk_mcu/p0_out [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4620_o,open_n38898}),
    .q({open_n38902,\u_cmsdk_mcu/p0_out [3]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4623|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n38903}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n38904}),
    .c({\u_cmsdk_mcu/p1_outen [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n105 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [3],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4623_o,open_n38921}),
    .q({open_n38925,\u_cmsdk_mcu/p1_altfunc [3]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~D*~(~B*~(~C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000011001110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4624|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b3/B1_0 ,open_n38926}),
    .b({_al_u4623_o,\u_cmsdk_mcu/p1_outen [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/p1_altfunc [3]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/p1_out [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4624_o,open_n38940}),
    .q({open_n38944,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [3]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"))
    \_al_u4627|_al_u4626  (
    .a({_al_u4624_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4625_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [3]}),
    .d({_al_u4626_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[3] }),
    .f({_al_u4627_o,_al_u4626_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~A*~(D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4629|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b3  (
    .a({_al_u4628_o,open_n38965}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .c({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .mi({open_n38977,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4629_o,_al_u4628_o}),
    .q({open_n38981,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [3]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~(~B*A)))"),
    //.LUT1("(D*~(C*~(~B*A)))"),
    .INIT_LUT0(16'b0010111100000000),
    .INIT_LUT1(16'b0010111100000000),
    .MODE("LOGIC"))
    \_al_u4630|_al_u4864  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o }),
    .b({_al_u4627_o,_al_u4861_o}),
    .c({_al_u4629_o,_al_u4863_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("((D@B)*(C@A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001001001001000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4631|_al_u5728  (
    .a({open_n39002,_al_u4106_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3],_al_u4141_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 }),
    .f({_al_u4631_o,_al_u5728_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0001011000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u4633|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b3_rom0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4633_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [3]}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*C)*~(B*A))"),
    //.LUTG0("~(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110101011000000),
    .INIT_LUTF1(16'b0000011101110111),
    .INIT_LUTG0(16'b1110101011000000),
    .INIT_LUTG1(16'b0000011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4634|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b3  (
    .a({\u_cmsdk_mcu/flash_hrdata [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4634_o,open_n39059}),
    .q({open_n39063,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [3]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    //.LUTF1("(A*~(D*C*B))"),
    //.LUTG0("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    //.LUTG1("(A*~(D*C*B))"),
    .INIT_LUTF0(16'b0001011000000000),
    .INIT_LUTF1(16'b0010101010101010),
    .INIT_LUTG0(16'b0001011000000000),
    .INIT_LUTG1(16'b0010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4636|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b3_rom0  (
    .a({_al_u4635_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}),
    .c({_al_u4580_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]}),
    .f({_al_u4636_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [3]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(D*~C*~B*~A)"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000000100000000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4637|_al_u4621  (
    .a({_al_u4621_o,_al_u4511_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [3],_al_u4618_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [3],_al_u4620_o}),
    .d({_al_u4636_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4637_o,_al_u4621_o}));
  // ../RTL/cortexm0ds_logic.v(17213)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4638|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,_al_u4638_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchiu6 }),
    .c({_al_u4637_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1839_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4638_o,open_n39129}),
    .q({open_n39133,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }));  // ../RTL/cortexm0ds_logic.v(17213)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u463|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b5  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({_al_u462_o,_al_u465_o}),
    .mi({open_n39139,\u_cmsdk_mcu/HADDR [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u463_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv }),
    .q({open_n39154,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[7] }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cortexm0ds_logic.v(18303)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010111000111111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4640|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6_reg  (
    .a({open_n39155,_al_u4500_o}),
    .b({_al_u4639_o,_al_u4501_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .mi({open_n39166,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchiu6 ,_al_u4639_o}),
    .q({open_n39171,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 }));  // ../RTL/cortexm0ds_logic.v(18303)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4642|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b4  (
    .a({_al_u1986_o,open_n39172}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39173}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n197 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4642_o,open_n39186}),
    .q({open_n39190,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [4]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4643|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n39191}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39192}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n242 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4643_o,open_n39209}),
    .q({open_n39213,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [4]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4645|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39214}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n39215}),
    .c({\u_cmsdk_mcu/p0_outen [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n62 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4645_o,open_n39228}),
    .q({open_n39232,\u_cmsdk_mcu/p0_outen [4]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4646|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b4  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [4]}),
    .b({_al_u4645_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [4],\u_cmsdk_mcu/p0_out [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4646_o,open_n39249}),
    .q({open_n39253,\u_cmsdk_mcu/p0_out [4]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4649|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39254}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n39255}),
    .c({\u_cmsdk_mcu/p1_outen [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n62 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4649_o,open_n39268}),
    .q({open_n39272,\u_cmsdk_mcu/p1_outen [4]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u464|_al_u472  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .d({_al_u463_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ,_al_u472_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~(~B*~(~C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011001110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4650|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b4/B1_0 ,open_n39299}),
    .b({_al_u4649_o,open_n39300}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/p1_outen [4]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/p1_out [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4650_o,open_n39314}),
    .q({open_n39318,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [4]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4651|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b4  (
    .a({_al_u1986_o,open_n39319}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39320}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n152 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [4],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4651_o,open_n39333}),
    .q({open_n39337,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [4]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4652|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n39338}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39339}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n279 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4652_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [4]}),
    .q({open_n39359,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[4] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~(~B*A)))"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(D*~(C*~(~B*A)))"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b0010111100000000),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0010111100000000),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4653|_al_u4656  (
    .a({_al_u4650_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o }),
    .b({_al_u4651_o,_al_u4653_o}),
    .c({_al_u1982_o,_al_u4655_o}),
    .d({_al_u4652_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]}),
    .f({_al_u4653_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [4]}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~A*~(D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4655|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b4  (
    .a({_al_u4654_o,open_n39384}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}),
    .c({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .mi({open_n39396,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4655_o,_al_u4654_o}),
    .q({open_n39400,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [4]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B@D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100000000110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4658|_al_u4850  (
    .b({open_n39403,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [3]}),
    .c({_al_u4605_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [4]}),
    .d({_al_u4657_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [2]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [4],_al_u4850_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B*~C*D+~A*B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1010011000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u4659|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b4_rom0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4659_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [4]}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110101011000000),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4660|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b4  (
    .a({\u_cmsdk_mcu/sram_hrdata [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4660_o,open_n39456}),
    .q({open_n39460,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [4]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(A*~(D*C*B))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(A*~(D*C*B))"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b0010101010101010),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b0010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4662|_al_u4661  (
    .a({_al_u4661_o,_al_u4659_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ,_al_u4660_o}),
    .c({_al_u4580_o,\u_cmsdk_mcu/flash_hrdata [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .f({_al_u4662_o,_al_u4661_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(D*~C*~B*~A)"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000000100000000),
    .MODE("LOGIC"))
    \_al_u4663|_al_u4647  (
    .a({_al_u4647_o,_al_u4511_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [4],_al_u4644_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [4],_al_u4646_o}),
    .d({_al_u4662_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4663_o,_al_u4647_o}));
  // ../RTL/cortexm0ds_logic.v(18706)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110100000001),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1100110100000001),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4664|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .c({_al_u4663_o,_al_u1841_o}),
    .clk(XTAL1_wire),
    .d({_al_u1841_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 }),
    .f({_al_u4664_o,open_n39523}),
    .q({open_n39527,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 }));  // ../RTL/cortexm0ds_logic.v(18706)
  // ../RTL/cortexm0ds_logic.v(17846)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4665|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,_al_u4664_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,_al_u4665_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tokax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4665_o,open_n39545}),
    .q({open_n39549,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgxpw6 }));  // ../RTL/cortexm0ds_logic.v(17846)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1010001100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4669|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b5_rom0  (
    .a({open_n39550,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4669_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [5]}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110101011000000),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4670|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b5  (
    .a({\u_cmsdk_mcu/sram_hrdata [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4670_o,open_n39583}),
    .q({open_n39587,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [5]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4672|_al_u4671  (
    .b({_al_u4671_o,\u_cmsdk_mcu/flash_hrdata [5]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({_al_u4669_o,_al_u4670_o}),
    .f({_al_u4672_o,_al_u4671_o}));
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001100000000),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1010001100000000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4673|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .b({_al_u4668_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}),
    .c({_al_u4672_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]}),
    .mi({open_n39617,\u_cmsdk_mcu/HADDR [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4673_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [5]}),
    .q({open_n39632,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_iop_gpio.v(387)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4675|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg3_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39633}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n39634}),
    .c({\u_cmsdk_mcu/p1_outen [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n88 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n109 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4675_o,open_n39651}),
    .q({open_n39655,\u_cmsdk_mcu/p1_altfunc [5]}));  // ../RTL/cmsdk_iop_gpio.v(387)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(~D*~(~B*~(~C*A)))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(~D*~(~B*~(~C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000000011001110),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000000011001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4676|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b5/B1_0 ,open_n39656}),
    .b({_al_u4675_o,\u_cmsdk_mcu/p1_outen [5]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/p1_altfunc [5]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/p1_out [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4676_o,open_n39674}),
    .q({open_n39678,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [5]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u4678|_al_u4677  (
    .a({open_n39679,_al_u1986_o}),
    .b({_al_u4676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4677_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [5]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [5]}),
    .f({_al_u4678_o,_al_u4677_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*B))"),
    //.LUTF1("(C*~B*~(~D*A))"),
    //.LUTG0("(~A*~(D*C*B))"),
    //.LUTG1("(C*~B*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b0011000000010000),
    .INIT_LUTG0(16'b0001010101010101),
    .INIT_LUTG1(16'b0011000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4681|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b5  (
    .a({_al_u1983_o,_al_u4669_o}),
    .b({_al_u4678_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .c({_al_u4679_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]}),
    .clk(XTAL1_wire),
    .d({_al_u4680_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]}),
    .mi({open_n39704,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4681_o,_al_u4679_o}),
    .q({open_n39719,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [5]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4682|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b5  (
    .a({_al_u1986_o,open_n39720}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39721}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n199 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4682_o,open_n39738}),
    .q({open_n39742,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [5]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000101111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4683|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n39743}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39744}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n244 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4683_o,open_n39757}),
    .q({open_n39761,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [5]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4685|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39762}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n39763}),
    .c({\u_cmsdk_mcu/p0_outen [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n64 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [5],\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4685_o,open_n39780}),
    .q({open_n39784,\u_cmsdk_mcu/p0_outen [5]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4686|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b5  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [5]}),
    .b({_al_u4685_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [5],\u_cmsdk_mcu/p0_out [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4686_o,open_n39801}),
    .q({open_n39805,\u_cmsdk_mcu/p0_out [5]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u4688|_al_u4687  (
    .a({_al_u4673_o,_al_u4511_o}),
    .b({_al_u4681_o,_al_u4684_o}),
    .c({_al_u4687_o,_al_u4686_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4688_o,_al_u4687_o}));
  // ../RTL/cortexm0ds_logic.v(18694)
  EG_PHY_LSLICE #(
    //.LUTF0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000100000001),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1111000100000001),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4689|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,_al_u1844_o}),
    .c({_al_u4688_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1844_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 }),
    .f({_al_u4689_o,open_n39844}),
    .q({open_n39848,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 }));  // ../RTL/cortexm0ds_logic.v(18694)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B*D))"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011110000),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u468|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b7  (
    .a({_al_u467_o,open_n39849}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n39860,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n26 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n285 }),
    .q({open_n39864,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [7]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cortexm0ds_logic.v(18699)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4690|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,_al_u4689_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,_al_u4690_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kakax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4690_o,open_n39878}),
    .q({open_n39882,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }));  // ../RTL/cortexm0ds_logic.v(18699)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4692|_al_u4515  (
    .a({_al_u1982_o,open_n39883}),
    .b({_al_u4515_o,open_n39884}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .d({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .f({_al_u4692_o,_al_u4515_o}));
  // ../RTL/cmsdk_iop_gpio.v(539)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000101111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4694|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg7_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n39909}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39910}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n283 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4694_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [6]}),
    .q({open_n39926,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[6] }));  // ../RTL/cmsdk_iop_gpio.v(539)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*~B*~(~D*A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*~B*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000001100000001),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000001100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4695|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b6  (
    .a({_al_u1983_o,open_n39927}),
    .b({_al_u4692_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]}),
    .c({_al_u4693_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({_al_u4694_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .mi({open_n39931,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4695_o,_al_u4693_o}),
    .q({open_n39946,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [6]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4697|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39947}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n39948}),
    .c({\u_cmsdk_mcu/p1_outen [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n66 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [6],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4697_o,open_n39961}),
    .q({open_n39965,\u_cmsdk_mcu/p1_outen [6]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~B*~(~C*A)))"),
    //.LUT1("(~D*~(~B*~(~C*A)))"),
    .INIT_LUT0(16'b0000000011001110),
    .INIT_LUT1(16'b0000000011001110),
    .MODE("LOGIC"))
    \_al_u4698|_al_u4833  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b6/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b8/B1_0 }),
    .b({_al_u4697_o,_al_u4832_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4698_o,_al_u4833_o}));
  // ../RTL/cmsdk_iop_gpio.v(425)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4699|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg4_b6  (
    .a({_al_u1986_o,open_n39986}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n39987}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n133 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n156 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [6],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4699_o,open_n40000}),
    .q({open_n40004,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [6]}));  // ../RTL/cmsdk_iop_gpio.v(425)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4701|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b6  (
    .a({_al_u1986_o,open_n40005}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40006}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n201 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [6],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4701_o,open_n40023}),
    .q({open_n40027,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [6]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4702|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n40028}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40029}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n246 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [6],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4702_o,open_n40046}),
    .q({open_n40050,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [6]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4704|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b6  (
    .a({open_n40051,\u_cmsdk_mcu/HWDATA [6]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/p0_out [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({_al_u4515_o,\u_cmsdk_mcu/p0_out [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4704_o,open_n40068}),
    .q({open_n40072,\u_cmsdk_mcu/p0_out [6]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4705|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40073}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n40074}),
    .c({\u_cmsdk_mcu/p0_outen [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n66 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [6],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4705_o,open_n40087}),
    .q({open_n40091,\u_cmsdk_mcu/p0_outen [6]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~(~C*~B)))"),
    //.LUTF1("(D*~(~C*~(B*~A)))"),
    //.LUTG0("(A*~(~D*~(~C*~B)))"),
    //.LUTG1("(D*~(~C*~(B*~A)))"),
    .INIT_LUTF0(16'b1010101000000010),
    .INIT_LUTF1(16'b1111010000000000),
    .INIT_LUTG0(16'b1010101000000010),
    .INIT_LUTG1(16'b1111010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4707|_al_u4706  (
    .a({_al_u4706_o,_al_u4703_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,_al_u4704_o}),
    .c({_al_u4692_o,_al_u4705_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [6],_al_u4706_o}));
  // ../RTL/cortexm0ds_logic.v(19867)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4708|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6_reg  (
    .a({\u_cmsdk_mcu/sram_hrdata [6],open_n40116}),
    .b({\u_cmsdk_mcu/flash_hrdata [6],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/flash_hrdata [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n40120,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4708_o,\u_cmsdk_mcu/u_ahb_rom/n13 [6]}),
    .q({open_n40135,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 }));  // ../RTL/cortexm0ds_logic.v(19867)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110101011000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1110101011000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4709|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b6  (
    .a({open_n40136,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({_al_u4708_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4709_o,open_n40153}),
    .q({open_n40157,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [6]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u470|_al_u467  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .d({_al_u467_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .f({_al_u470_o,_al_u467_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D+~A*B*C*D)"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D+~A*B*C*D)"),
    //.LUTG1("(D*C*~B*A)"),
    .INIT_LUTF0(16'b0101000100010000),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0101000100010000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4710|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b2_rom0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b6_sel_is_13_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u4711|_al_u4668  (
    .b({_al_u4709_o,open_n40212}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b6_sel_is_13_o ,_al_u4580_o}),
    .d({_al_u4668_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o }),
    .f({_al_u4711_o,_al_u4668_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(C*~B*~(D*~A))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(C*~B*~(D*~A))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0010000000110000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0010000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4712|_al_u4700  (
    .a({_al_u4700_o,_al_u4695_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o }),
    .c({_al_u4711_o,_al_u4698_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],_al_u4699_o}),
    .f({_al_u4712_o,_al_u4700_o}));
  // ../RTL/cortexm0ds_logic.v(18693)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110100000001),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1100110100000001),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4713|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .c({_al_u4712_o,_al_u1846_o}),
    .clk(XTAL1_wire),
    .d({_al_u1846_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 }),
    .f({_al_u4713_o,open_n40275}),
    .q({open_n40279,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 }));  // ../RTL/cortexm0ds_logic.v(18693)
  // ../RTL/cortexm0ds_logic.v(18632)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4714|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,_al_u4713_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5hiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8kax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5hiu6 ,open_n40297}),
    .q({open_n40301,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }));  // ../RTL/cortexm0ds_logic.v(18632)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1010001000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1010001000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4716|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b7_rom0  (
    .a({open_n40302,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4716_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [7]}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*C)*~(B*A))"),
    //.LUTG0("~(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110101011000000),
    .INIT_LUTF1(16'b0000011101110111),
    .INIT_LUTG0(16'b1110101011000000),
    .INIT_LUTG1(16'b0000011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4717|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b7  (
    .a({\u_cmsdk_mcu/sram_hrdata [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4717_o,open_n40343}),
    .q({open_n40347,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [7]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u4719|_al_u4718  (
    .b({_al_u4718_o,\u_cmsdk_mcu/flash_hrdata [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}),
    .d({_al_u4716_o,_al_u4717_o}),
    .f({_al_u4719_o,_al_u4718_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u471|_al_u458  (
    .c({_al_u470_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u4720|_al_u4796  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [5],open_n40398}),
    .b({_al_u4668_o,_al_u4795_o}),
    .c({_al_u4719_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [7],_al_u4787_o}),
    .f({_al_u4720_o,_al_u4796_o}));
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4722|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40419}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n40420}),
    .c({\u_cmsdk_mcu/p1_outen [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n68 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4722_o,open_n40433}),
    .q({open_n40437,\u_cmsdk_mcu/p1_outen [7]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~(~B*~(~C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011001110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4723|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b7/B1_0 ,open_n40438}),
    .b({_al_u4722_o,open_n40439}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/p1_outen [7]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/p1_out [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4723_o,open_n40453}),
    .q({open_n40457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [7]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4724|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg5_b7  (
    .a({_al_u1986_o,open_n40458}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40459}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n203 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4724_o,open_n40476}),
    .q({open_n40480,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [7]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~(~D*A))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b0000001100000001),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u4725|_al_u4589  (
    .a({open_n40481,_al_u1983_o}),
    .b({_al_u4723_o,_al_u4586_o}),
    .c({_al_u4724_o,_al_u4587_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,_al_u4588_o}),
    .f({_al_u4725_o,_al_u4589_o}));
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000101111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4727|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg6_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n40502}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40503}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n248 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[7] ,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4727_o,open_n40516}),
    .q({open_n40520,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [7]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*B))"),
    //.LUTF1("(C*~B*~(~D*A))"),
    //.LUTG0("(~A*~(D*C*B))"),
    //.LUTG1("(C*~B*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b0011000000010000),
    .INIT_LUTG0(16'b0001010101010101),
    .INIT_LUTG1(16'b0011000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4728|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b7  (
    .a({_al_u1983_o,_al_u4716_o}),
    .b({_al_u4725_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .c({_al_u4726_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}),
    .clk(XTAL1_wire),
    .d({_al_u4727_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]}),
    .mi({open_n40525,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4728_o,_al_u4726_o}),
    .q({open_n40540,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [7]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(463)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4729|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg5_b7  (
    .a({_al_u1986_o,open_n40541}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40542}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n178 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n203 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4729_o,open_n40559}),
    .q({open_n40563,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [7]}));  // ../RTL/cmsdk_iop_gpio.v(463)
  // ../RTL/cmsdk_iop_gpio.v(501)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4730|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg6_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n40564}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40565}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n223 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n248 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4730_o,open_n40582}),
    .q({open_n40586,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [7]}));  // ../RTL/cmsdk_iop_gpio.v(501)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4732|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg2_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40587}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n40588}),
    .c({\u_cmsdk_mcu/p0_outen [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n68 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_altfunc [7],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4732_o,open_n40605}),
    .q({open_n40609,\u_cmsdk_mcu/p0_outen [7]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4733|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b7  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [7]}),
    .b({_al_u4732_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [7],\u_cmsdk_mcu/p0_out [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4733_o,open_n40626}),
    .q({open_n40630,\u_cmsdk_mcu/p0_out [7]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4735|_al_u4734  (
    .a({_al_u4720_o,_al_u4511_o}),
    .b({_al_u4728_o,_al_u4731_o}),
    .c({_al_u4734_o,_al_u4733_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4735_o,_al_u4734_o}));
  // ../RTL/cortexm0ds_logic.v(18690)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4736|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,_al_u4736_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2hiu6 }),
    .c({_al_u4735_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1848_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4736_o,open_n40668}),
    .q({open_n40672,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }));  // ../RTL/cortexm0ds_logic.v(18690)
  // ../RTL/cortexm0ds_logic.v(18304)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010111000111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0010111000111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4738|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6_reg  (
    .a({open_n40673,_al_u4500_o}),
    .b({_al_u4737_o,_al_u4501_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .mi({open_n40677,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2hiu6 ,_al_u4737_o}),
    .q({open_n40693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 }));  // ../RTL/cortexm0ds_logic.v(18304)
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u473|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b0  (
    .a({open_n40694,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }),
    .b({open_n40695,_al_u472_o}),
    .c({_al_u472_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({_al_u463_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .mi({open_n40706,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 }),
    .q({open_n40710,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]}));  // ../RTL/gpio_apbif.v(262)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"))
    \_al_u4740|_al_u4890  (
    .a({_al_u1986_o,_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [15]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [15]}),
    .f({_al_u4740_o,_al_u4890_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4742|_al_u4741  (
    .a({open_n40731,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4741_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [9]}),
    .d({_al_u4740_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [9]}),
    .f({_al_u4742_o,_al_u4741_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1100100001000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1100100001000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4743|_al_u4893  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c({\u_cmsdk_mcu/p0_outen [9],\u_cmsdk_mcu/p0_outen [15]}),
    .d({\u_cmsdk_mcu/p0_altfunc [9],\u_cmsdk_mcu/p0_altfunc [15]}),
    .f({_al_u4743_o,_al_u4893_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4744|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b9  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [9]}),
    .b({_al_u4743_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4:3]),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [9],\u_cmsdk_mcu/p0_out [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4744_o,open_n40792}),
    .q({open_n40796,\u_cmsdk_mcu/p0_out [9]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4746|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b9  (
    .a({\u_cmsdk_mcu/sram_hrdata [9],open_n40797}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],open_n40798}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4746_o,open_n40811}),
    .q({open_n40815,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [9]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4747|_al_u4745  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [9],_al_u4511_o}),
    .b({_al_u4746_o,_al_u4742_o}),
    .c({\u_cmsdk_mcu/flash_hrdata [9],_al_u4744_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4747_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [9]}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4749|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b9  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n40840}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n40841}),
    .c({\u_cmsdk_mcu/p1_outen [9],\u_cmsdk_mcu/p1_outen [9]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [9],\u_cmsdk_mcu/p1_out [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4749_o,open_n40859}),
    .q({open_n40863,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [9]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~B*~(~C*A)))"),
    //.LUT1("(~D*~(~B*~(~C*A)))"),
    .INIT_LUT0(16'b0000000011001110),
    .INIT_LUT1(16'b0000000011001110),
    .MODE("LOGIC"))
    \_al_u4750|_al_u4802  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b9/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b12/B1_0 }),
    .b({_al_u4749_o,_al_u4801_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4750_o,_al_u4802_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4752|_al_u4751  (
    .a({open_n40884,_al_u1986_o}),
    .b({_al_u4750_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4751_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [9]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [9]}),
    .f({_al_u4752_o,_al_u4751_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4755|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b9  (
    .a({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4752_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4753_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .clk(XTAL1_wire),
    .d({_al_u4754_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]}),
    .mi({open_n40920,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4755_o,_al_u4753_o}),
    .q({open_n40924,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [9]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(D*~B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(C*~A*~(D*~B))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b0100000001010000),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4756|_al_u4529  (
    .a({open_n40925,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [14]}),
    .b({_al_u4755_o,_al_u4526_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],_al_u4528_o}),
    .d({_al_u4747_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]}),
    .f({_al_u4756_o,_al_u4529_o}));
  // ../RTL/cortexm0ds_logic.v(18671)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110100000001),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4757|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .c({_al_u4756_o,_al_u1852_o}),
    .clk(XTAL1_wire),
    .d({_al_u1852_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 }),
    .f({_al_u4757_o,open_n40964}),
    .q({open_n40968,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 }));  // ../RTL/cortexm0ds_logic.v(18671)
  // ../RTL/cortexm0ds_logic.v(18676)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4758|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,_al_u4757_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,_al_u4758_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sujax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4758_o,open_n40986}),
    .q({open_n40990,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }));  // ../RTL/cortexm0ds_logic.v(18676)
  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u475|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5]}),
    .b({_al_u473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [5]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b5/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .mi({open_n41001,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u475_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b5/B1_0 }),
    .q({open_n41005,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [5]}));  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"))
    \_al_u4760|_al_u4878  (
    .a({_al_u1986_o,_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [13]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [13]}),
    .f({_al_u4760_o,_al_u4878_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4762|_al_u4761  (
    .a({open_n41026,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4761_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [10]}),
    .d({_al_u4760_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [10]}),
    .f({_al_u4762_o,_al_u4761_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1100100001000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1100100001000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4763|_al_u4881  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c({\u_cmsdk_mcu/p0_outen [10],\u_cmsdk_mcu/p0_outen [13]}),
    .d({\u_cmsdk_mcu/p0_altfunc [10],\u_cmsdk_mcu/p0_altfunc [13]}),
    .f({_al_u4763_o,_al_u4881_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b0011000100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4764|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b10  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [10]}),
    .b({_al_u4763_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [10],\u_cmsdk_mcu/p0_out [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4764_o,open_n41083}),
    .q({open_n41087,\u_cmsdk_mcu/p0_out [10]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*C)*~(B*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000011101110111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4766|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b10  (
    .a({\u_cmsdk_mcu/sram_hrdata [10],open_n41088}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],open_n41089}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [10]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4766_o,open_n41106}),
    .q({open_n41110,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [10]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u4767|_al_u4765  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [10],_al_u4511_o}),
    .b({_al_u4766_o,_al_u4762_o}),
    .c({\u_cmsdk_mcu/flash_hrdata [10],_al_u4764_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4767_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [10]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4770|_al_u4769  (
    .a({open_n41131,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4769_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [10]}),
    .d({_al_u4768_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[10] }),
    .f({_al_u4770_o,_al_u4769_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4772|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b10  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n41156}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n41157}),
    .c({\u_cmsdk_mcu/p1_outen [10],\u_cmsdk_mcu/p1_outen [10]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [10],\u_cmsdk_mcu/p1_out [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4772_o,open_n41175}),
    .q({open_n41179,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [10]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~B*~(~C*A)))"),
    //.LUTF1("(~D*~(~B*~(~C*A)))"),
    //.LUTG0("(~D*~(~B*~(~C*A)))"),
    //.LUTG1("(~D*~(~B*~(~C*A)))"),
    .INIT_LUTF0(16'b0000000011001110),
    .INIT_LUTF1(16'b0000000011001110),
    .INIT_LUTG0(16'b0000000011001110),
    .INIT_LUTG1(16'b0000000011001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4773|_al_u4793  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b10/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b11/B1_0 }),
    .b({_al_u4772_o,_al_u4792_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4773_o,_al_u4793_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*~A)"),
    //.LUTF1("(~D*~(A*~(~C*B)))"),
    //.LUTG0("(D*C*B*~A)"),
    //.LUTG1("(~D*~(A*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000000000000),
    .INIT_LUTF1(16'b0000000001011101),
    .INIT_LUTG0(16'b0100000000000000),
    .INIT_LUTG1(16'b0000000001011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4775|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b10  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4770_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4773_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .clk(XTAL1_wire),
    .d({_al_u4774_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]}),
    .mi({open_n41208,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4775_o,_al_u4774_o}),
    .q({open_n41223,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [10]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u4776|_al_u4836  (
    .b({_al_u4775_o,_al_u4835_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]}),
    .d({_al_u4767_o,_al_u4827_o}),
    .f({_al_u4776_o,_al_u4836_o}));
  // ../RTL/cortexm0ds_logic.v(18664)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110100000001),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1100110100000001),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4777|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .c({_al_u4776_o,_al_u1854_o}),
    .clk(XTAL1_wire),
    .d({_al_u1854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 }),
    .f({_al_u4777_o,open_n41264}),
    .q({open_n41268,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 }));  // ../RTL/cortexm0ds_logic.v(18664)
  // ../RTL/cortexm0ds_logic.v(18669)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4778|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,_al_u4777_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epciu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqjax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Epciu6 ,open_n41282}),
    .q({open_n41286,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }));  // ../RTL/cortexm0ds_logic.v(18669)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4780|_al_u4844  (
    .a({_al_u1986_o,_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [0]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [0]}),
    .f({_al_u4780_o,_al_u4844_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4782|_al_u4781  (
    .a({open_n41311,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4781_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [11]}),
    .d({_al_u4780_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [11]}),
    .f({_al_u4782_o,_al_u4781_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b1100100001000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"))
    \_al_u4783|_al_u4847  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c({\u_cmsdk_mcu/p0_outen [11],\u_cmsdk_mcu/p0_outen [0]}),
    .d({\u_cmsdk_mcu/p0_altfunc [11],\u_cmsdk_mcu/p0_altfunc [0]}),
    .f({_al_u4783_o,_al_u4847_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4784|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b11  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [11]}),
    .b({_al_u4783_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [11],\u_cmsdk_mcu/p0_out [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4784_o,open_n41372}),
    .q({open_n41376,\u_cmsdk_mcu/p0_out [11]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4787|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b11  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [11],open_n41377}),
    .b({_al_u4786_o,open_n41378}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [11]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4787_o,open_n41395}),
    .q({open_n41399,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [11]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u478|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [4]}),
    .b({_al_u473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [4]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b4/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .mi({open_n41403,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b4/B1_0 }),
    .q({open_n41418,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [4]}));  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4790|_al_u4789  (
    .a({open_n41419,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4789_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [11]}),
    .d({_al_u4788_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[11] }),
    .f({_al_u4790_o,_al_u4789_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4792|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b11  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n41440}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n41441}),
    .c({\u_cmsdk_mcu/p1_outen [11],\u_cmsdk_mcu/p1_outen [11]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [11],\u_cmsdk_mcu/p1_out [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4792_o,open_n41455}),
    .q({open_n41459,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [11]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*~A)"),
    //.LUTF1("(~D*~(A*~(~C*B)))"),
    //.LUTG0("(D*C*B*~A)"),
    //.LUTG1("(~D*~(A*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000000000000),
    .INIT_LUTF1(16'b0000000001011101),
    .INIT_LUTG0(16'b0100000000000000),
    .INIT_LUTG1(16'b0000000001011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4795|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b11  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4790_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4793_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .clk(XTAL1_wire),
    .d({_al_u4794_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]}),
    .mi({open_n41464,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4795_o,_al_u4794_o}),
    .q({open_n41479,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [11]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cortexm0ds_logic.v(18657)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110100000001),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1100110100000001),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4797|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .c({_al_u4796_o,_al_u1856_o}),
    .clk(XTAL1_wire),
    .d({_al_u1856_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 }),
    .f({_al_u4797_o,open_n41498}),
    .q({open_n41502,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 }));  // ../RTL/cortexm0ds_logic.v(18657)
  // ../RTL/cortexm0ds_logic.v(18662)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4798|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,_al_u4797_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anciu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smjax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Anciu6 ,open_n41516}),
    .q({open_n41520,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }));  // ../RTL/cortexm0ds_logic.v(18662)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4801|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b12  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n41521}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n41522}),
    .c({\u_cmsdk_mcu/p1_outen [12],\u_cmsdk_mcu/p1_outen [12]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [12],\u_cmsdk_mcu/p1_out [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4801_o,open_n41536}),
    .q({open_n41540,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [12]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u4804|_al_u4803  (
    .a({open_n41541,_al_u1986_o}),
    .b({_al_u4802_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4803_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [12]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [12]}),
    .f({_al_u4804_o,_al_u4803_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4807|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b12  (
    .a({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4804_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4805_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}),
    .clk(XTAL1_wire),
    .d({_al_u4806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]}),
    .mi({open_n41573,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4807_o,_al_u4805_o}),
    .q({open_n41577,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [12]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4808|_al_u4820  (
    .a({_al_u1986_o,_al_u1986_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inten_padded [8]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_inttype_padded [8]}),
    .f({_al_u4808_o,_al_u4820_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4810|_al_u4809  (
    .a({open_n41602,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4809_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [12]}),
    .d({_al_u4808_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [12]}),
    .f({_al_u4810_o,_al_u4809_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b1100100001000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"))
    \_al_u4811|_al_u4823  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c({\u_cmsdk_mcu/p0_outen [12],\u_cmsdk_mcu/p0_outen [8]}),
    .d({\u_cmsdk_mcu/p0_altfunc [12],\u_cmsdk_mcu/p0_altfunc [8]}),
    .f({_al_u4811_o,_al_u4823_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b0011000100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4812|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b12  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [12]}),
    .b({_al_u4811_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [12],\u_cmsdk_mcu/p0_out [12]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4812_o,open_n41659}),
    .q({open_n41663,\u_cmsdk_mcu/p0_out [12]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4815|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b12  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n41664}),
    .b({_al_u4814_o,open_n41665}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [12]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4815_o,open_n41678}),
    .q({open_n41682,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [12]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(C*~B*~(D*~A))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(C*~B*~(D*~A))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0010000000110000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0010000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4816|_al_u4813  (
    .a({_al_u4807_o,_al_u4511_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [12],_al_u4810_o}),
    .c({_al_u4815_o,_al_u4812_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4816_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [12]}));
  // ../RTL/cortexm0ds_logic.v(18650)
  EG_PHY_MSLICE #(
    //.LUT0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100000001),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4817|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,_al_u1859_o}),
    .c({_al_u4816_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1859_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 }),
    .f({_al_u4817_o,open_n41721}),
    .q({open_n41725,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 }));  // ../RTL/cortexm0ds_logic.v(18650)
  // ../RTL/cortexm0ds_logic.v(18655)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4818|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,_al_u4817_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkciu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sijax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkciu6 ,open_n41739}),
    .q({open_n41743,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Skjax6 }));  // ../RTL/cortexm0ds_logic.v(18655)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4822|_al_u4821  (
    .a({open_n41744,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4821_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [8]}),
    .d({_al_u4820_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [8]}),
    .f({_al_u4822_o,_al_u4821_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4824|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b8  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [8]}),
    .b({_al_u4823_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [8],\u_cmsdk_mcu/p0_out [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4824_o,open_n41781}),
    .q({open_n41785,\u_cmsdk_mcu/p0_out [8]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4827|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b8  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [8],open_n41786}),
    .b({_al_u4826_o,open_n41787}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4827_o,open_n41800}),
    .q({open_n41804,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [8]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~D*A*~(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0000000010101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u482|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [3]}),
    .b({_al_u480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [3]}),
    .c({_al_u481_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .mi({open_n41815,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u482_o,_al_u481_o}),
    .q({open_n41819,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [3]}));  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4830|_al_u4829  (
    .a({open_n41820,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4829_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [8]}),
    .d({_al_u4828_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[8] }),
    .f({_al_u4830_o,_al_u4829_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4832|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b8  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n41845}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n41846}),
    .c({\u_cmsdk_mcu/p1_outen [8],\u_cmsdk_mcu/p1_outen [8]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [8],\u_cmsdk_mcu/p1_out [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4832_o,open_n41864}),
    .q({open_n41868,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [8]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~D*~(A*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000000001011101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4835|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b8  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4830_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4833_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .clk(XTAL1_wire),
    .d({_al_u4834_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]}),
    .mi({open_n41880,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4835_o,_al_u4834_o}),
    .q({open_n41884,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [8]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cortexm0ds_logic.v(18678)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110100000001),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1100110100000001),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4837|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .c({_al_u4836_o,_al_u1850_o}),
    .clk(XTAL1_wire),
    .d({_al_u1850_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 }),
    .f({_al_u4837_o,open_n41903}),
    .q({open_n41907,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 }));  // ../RTL/cortexm0ds_logic.v(18678)
  // ../RTL/cortexm0ds_logic.v(18683)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4838|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,_al_u4837_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,_al_u4838_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4838_o,open_n41921}),
    .q({open_n41925,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }));  // ../RTL/cortexm0ds_logic.v(18683)
  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u483|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b3  (
    .b({_al_u482_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ,_al_u483_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u483_o,open_n41940}),
    .q({open_n41944,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [3]}));  // ../RTL/cmsdk_apb_uart.v(303)
  // ../RTL/cmsdk_mcu_sysctrl.v(290)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4840|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2],_al_u497_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3],_al_u499_o}),
    .c({\u_cmsdk_mcu/LOCKUPRESET ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_write ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/remap_ctrl ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}),
    .mi({open_n41955,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux3_b0/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_lockupreset_write }),
    .q({open_n41959,\u_cmsdk_mcu/LOCKUPRESET }));  // ../RTL/cmsdk_mcu_sysctrl.v(290)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*A)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(D*~C*~B*A)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4841|_al_u2993  (
    .a({open_n41960,_al_u2992_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux3_b0/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4:3]),
    .d({_al_u2992_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}),
    .f({_al_u4841_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*A*~(D*~B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*A*~(D*~B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000100000001010),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4842|_al_u4581  (
    .a({open_n41985,_al_u4568_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux6_b3_sel_is_2_o ,_al_u4571_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [1]}),
    .d({_al_u4841_o,_al_u4580_o}),
    .f({_al_u4842_o,_al_u4581_o}));
  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*A)))"),
    //.LUTF1("(C*~(A*~(D*B)))"),
    //.LUTG0("~(~D*~(C*~(B*A)))"),
    //.LUTG1("(C*~(A*~(D*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111101110000),
    .INIT_LUTF1(16'b1101000001010000),
    .INIT_LUTG0(16'b1111111101110000),
    .INIT_LUTG1(16'b1101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4843|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg2_b0  (
    .a({_al_u4842_o,\u_cmsdk_mcu/HWDATA [0]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n34_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_write }),
    .c({_al_u4580_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo_en ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [0],\u_cmsdk_mcu/SYSRESETREQ }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n35 [0],open_n42026}),
    .q({open_n42030,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_resetinfo [0]}));  // ../RTL/cmsdk_mcu_sysctrl.v(318)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4846|_al_u4845  (
    .a({open_n42031,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4845_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [0]}),
    .d({_al_u4844_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [0]}),
    .f({_al_u4846_o,_al_u4845_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b0011000100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4848|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b0  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [0]}),
    .b({_al_u4847_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [0],\u_cmsdk_mcu/p0_out [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4848_o,open_n42068}),
    .q({open_n42072,\u_cmsdk_mcu/p0_out [0]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u4851|_al_u4855  (
    .a({_al_u4657_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [2]}),
    .b({_al_u4850_o,_al_u4851_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [1],_al_u4854_o}),
    .f({_al_u4851_o,_al_u4855_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1101010000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1101010000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4852|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux2_b0_rom0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4852_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [0]}));
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110101011000000),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4853|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b0  (
    .a({\u_cmsdk_mcu/flash_hrdata [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4853_o,open_n42129}),
    .q({open_n42133,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [0]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u4854|_al_u2009  (
    .a({_al_u4852_o,open_n42134}),
    .b({_al_u4853_o,\u_cmsdk_mcu/sram_hrdata [0]}),
    .c({\u_cmsdk_mcu/sram_hrdata [0],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1],\u_cmsdk_mcu/HWDATA [0]}),
    .f({_al_u4854_o,\u_cmsdk_mcu/u_ahb_ram/n13 [0]}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011001000010000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011001000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4856|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],open_n42155}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n42156}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0],\u_cmsdk_mcu/p1_outen [0]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [0],\u_cmsdk_mcu/p1_out [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b0/B1_0 ,open_n42174}),
    .q({open_n42178,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [0]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(348)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4857|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg2_b0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n42179}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n42180}),
    .c({\u_cmsdk_mcu/p1_outen [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n43 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n54 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [0],\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4857_o,open_n42193}),
    .q({open_n42197,\u_cmsdk_mcu/p1_outen [0]}));  // ../RTL/cmsdk_iop_gpio.v(348)
  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(~C*~(B*D))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111110011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u485|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b4  (
    .b({open_n42200,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [4],\u_cmsdk_mcu/HWDATA [4]}),
    .mi({open_n42204,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n279 }),
    .q({open_n42219,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [4]}));  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4861|_al_u4860  (
    .a({_al_u4858_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u4859_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [0]}),
    .d({_al_u4860_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[0] }),
    .f({_al_u4861_o,_al_u4860_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~A*~(D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4863|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b0  (
    .a({_al_u4862_o,open_n42244}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .c({_al_u4566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n13 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .mi({open_n42249,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4863_o,_al_u4862_o}),
    .q({open_n42264,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [0]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(~D*C*~B*~A)"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000000000010000),
    .MODE("LOGIC"))
    \_al_u4865|_al_u4849  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n35 [0],_al_u4511_o}),
    .b({_al_u4849_o,_al_u4846_o}),
    .c({_al_u4855_o,_al_u4848_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n33 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4865_o,_al_u4849_o}));
  // ../RTL/cortexm0ds_logic.v(17655)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4866|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,_al_u4866_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3biu6 }),
    .c({_al_u4865_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4866_o,open_n42298}),
    .q({open_n42302,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }));  // ../RTL/cortexm0ds_logic.v(17655)
  // ../RTL/cortexm0ds_logic.v(18177)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010111000111111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0010111000111111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4868|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6_reg  (
    .a({open_n42303,_al_u4500_o}),
    .b({_al_u4867_o,_al_u4501_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .mi({open_n42307,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3biu6 ,_al_u4867_o}),
    .q({open_n42323,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 }));  // ../RTL/cortexm0ds_logic.v(18177)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4871|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b13  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],open_n42324}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],open_n42325}),
    .c({\u_cmsdk_mcu/p1_outen [13],\u_cmsdk_mcu/p1_outen [13]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_altfunc [13],\u_cmsdk_mcu/p1_out [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4871_o,open_n42343}),
    .q({open_n42347,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [13]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u4874|_al_u4873  (
    .a({open_n42348,_al_u1986_o}),
    .b({_al_u4872_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4873_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [13]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [13]}),
    .f({_al_u4874_o,_al_u4873_o}));
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4877|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b13  (
    .a({_al_u1983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4874_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4875_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]}),
    .clk(XTAL1_wire),
    .d({_al_u4876_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]}),
    .mi({open_n42380,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4877_o,_al_u4875_o}),
    .q({open_n42384,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [13]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*D))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("~(~C*~(B*D))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011110000),
    .INIT_LUTF1(16'b1111010100111111),
    .INIT_LUTG0(16'b1111110011110000),
    .INIT_LUTG1(16'b1111010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u487|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [2],open_n42385}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_overrun ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [2]}),
    .mi({open_n42389,\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u487_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n275 }),
    .q({open_n42404,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [2]}));  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1000101111001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4880|_al_u4879  (
    .a({open_n42405,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4879_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [13]}),
    .d({_al_u4878_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [13]}),
    .f({_al_u4880_o,_al_u4879_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b0011000100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4882|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b13  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [13]}),
    .b({_al_u4881_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [13],\u_cmsdk_mcu/p0_out [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4882_o,open_n42438}),
    .q({open_n42442,\u_cmsdk_mcu/p0_out [13]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4885|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b13  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n42443}),
    .b({_al_u4884_o,open_n42444}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [13]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4885_o,open_n42457}),
    .q({open_n42461,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [13]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(C*~B*~(D*~A))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0010000000110000),
    .MODE("LOGIC"))
    \_al_u4886|_al_u4883  (
    .a({_al_u4877_o,_al_u4511_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [13],_al_u4880_o}),
    .c({_al_u4885_o,_al_u4882_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4886_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [13]}));
  // ../RTL/cortexm0ds_logic.v(18649)
  EG_PHY_MSLICE #(
    //.LUT0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100000001),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4887|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pp7iu6 ,_al_u1862_o}),
    .c({_al_u4886_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({_al_u1862_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 }),
    .f({_al_u4887_o,open_n42496}),
    .q({open_n42500,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 }));  // ../RTL/cortexm0ds_logic.v(18649)
  // ../RTL/cortexm0ds_logic.v(18060)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4888|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,_al_u4887_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U28iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sgjax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U28iu6 ,open_n42514}),
    .q({open_n42518,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }));  // ../RTL/cortexm0ds_logic.v(18060)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(~D*A*~(C*B))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b0000000000101010),
    .MODE("LOGIC"))
    \_al_u488|_al_u486  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/uart0_txovrint }),
    .b({_al_u486_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [2]}),
    .c({_al_u487_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .f({_al_u488_o,_al_u486_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1000101111001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1000101111001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4892|_al_u4891  (
    .a({open_n42539,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4891_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intpol_padded [15]}),
    .d({_al_u4890_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_intr [15]}),
    .f({_al_u4892_o,_al_u4891_o}));
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4894|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg1_b15  (
    .a({_al_u4515_o,\u_cmsdk_mcu/HWDATA [15]}),
    .b({_al_u4893_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p0_out [15],\u_cmsdk_mcu/p0_out [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4894_o,open_n42580}),
    .q({open_n42584,\u_cmsdk_mcu/p0_out [15]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTF1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG1("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010010110100001),
    .INIT_LUTF1(16'b1000101111001111),
    .INIT_LUTG0(16'b0010010110100001),
    .INIT_LUTG1(16'b1000101111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4897|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg8_b15  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intpol_padded [15]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n304 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/GPIOINT[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [15]}),
    .mi({open_n42588,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4897_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_raw_int [15]}),
    .q({open_n42603,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_last_datain [15]}));  // ../RTL/cmsdk_iop_gpio.v(561)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4898|_al_u4896  (
    .a({open_n42604,_al_u1986_o}),
    .b({_al_u1982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({_al_u4897_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inten_padded [15]}),
    .d({_al_u4896_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_inttype_padded [15]}),
    .f({_al_u4898_o,_al_u4896_o}));
  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u489|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b2  (
    .b({_al_u488_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ,_al_u489_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u489_o,open_n42639}),
    .q({open_n42643,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [2]}));  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(~B*~(~C*A)))"),
    .INIT_LUT0(16'b1100100001000000),
    .INIT_LUT1(16'b0000000011001110),
    .MODE("LOGIC"))
    \_al_u4901|_al_u4900  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b15/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .b({_al_u4900_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4],\u_cmsdk_mcu/p1_outen [15]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/p1_altfunc [15]}),
    .f({_al_u4901_o,_al_u4900_o}));
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*~A)"),
    //.LUTF1("(~D*~(A*~(~C*B)))"),
    //.LUTG0("(D*C*B*~A)"),
    //.LUTG1("(~D*~(A*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000000000000),
    .INIT_LUTF1(16'b0000000001011101),
    .INIT_LUTG0(16'b0100000000000000),
    .INIT_LUTG1(16'b0000000001011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4903|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b9  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/mux4_b10_sel_is_4_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .b({_al_u4898_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .c({_al_u4901_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}),
    .clk(XTAL1_wire),
    .d({_al_u4902_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]}),
    .mi({open_n42668,\u_cmsdk_mcu/HADDR [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4903_o,_al_u4902_o}),
    .q({open_n42683,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4905|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg3_b15  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n37 [14],open_n42684}),
    .b({_al_u4904_o,open_n42685}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [15]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4905_o,open_n42702}),
    .q({open_n42706,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/rwdata_reg [15]}));  // ../RTL/cmsdk_ahb_to_apb.v(265)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(C*~A*~(D*~B))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(C*~A*~(D*~B))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0100000001010000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0100000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4906|_al_u4895  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [15],_al_u4511_o}),
    .b({_al_u4903_o,_al_u4892_o}),
    .c({_al_u4905_o,_al_u4894_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .f({_al_u4906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n31 [15]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0100010111001111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u4907|_al_u6834  (
    .a({open_n42731,_al_u6087_o}),
    .b({open_n42732,_al_u4906_o}),
    .c({_al_u4533_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({_al_u4906_o,_al_u6817_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 }));
  // ../RTL/cortexm0ds_logic.v(18648)
  EG_PHY_LSLICE #(
    //.LUTF0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000100000001),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000100000001),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4908|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M15iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uy4iu6 ,_al_u1865_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 }),
    .f({_al_u4908_o,open_n42771}),
    .q({open_n42775,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sejax6 }));  // ../RTL/cortexm0ds_logic.v(18648)
  // ../RTL/cortexm0ds_logic.v(17876)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(~C*B))"),
    //.LUT1("(C*A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011111111),
    .INIT_LUT1(16'b0010000010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4910|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6_reg  (
    .a({_al_u4908_o,open_n42776}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kq7iu6 }),
    .c({_al_u4909_o,_al_u1865_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 ,_al_u4910_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4910_o,open_n42790}),
    .q({open_n42794,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }));  // ../RTL/cortexm0ds_logic.v(17876)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4913|_al_u4912  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv }),
    .d({_al_u4912_o,_al_u4368_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ,_al_u4912_o}));
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~((D*~C))*~(A)+B*(D*~C)*~(A)+~(B)*(D*~C)*A+B*(D*~C)*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~((D*~C))*~(A)+B*(D*~C)*~(A)+~(B)*(D*~C)*A+B*(D*~C)*A)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100111001000100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0100111001000100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4914|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b0  (
    .a({open_n42823,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .b({open_n42824,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ,_al_u4914_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4914_o,\u_cmsdk_mcu/HADDR [0]}),
    .q({open_n42845,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [0]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4917|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b0  (
    .b({_al_u4548_o,_al_u4552_o}),
    .c({_al_u4553_o,_al_u4553_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({_al_u4916_o,_al_u4548_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4917_o,\u_cmsdk_mcu/flash_hsel }),
    .q({open_n42867,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [0]}));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*~(~C*~A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111101011001000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4919|_al_u5798  (
    .a({open_n42868,_al_u4061_o}),
    .b({_al_u4061_o,_al_u4126_o}),
    .c({_al_u4066_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 }),
    .d({_al_u4918_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 }),
    .f({_al_u4919_o,_al_u5798_o}));
  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000101000001100),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000101000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u491|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b0  (
    .a({uart0_txen_pad,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [0],_al_u370_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]}),
    .mi({open_n42892,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u491_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample }),
    .q({open_n42907,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [0]}));  // ../RTL/cmsdk_apb_uart.v(603)
  // ../RTL/cortexm0ds_logic.v(18042)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4920|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6_reg  (
    .a({open_n42908,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [7]}),
    .mi({open_n42912,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 }),
    .f({_al_u4920_o,_al_u5824_o}),
    .q({open_n42928,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 }));  // ../RTL/cortexm0ds_logic.v(18042)
  // ../RTL/cortexm0ds_logic.v(19993)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4922|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6_reg  (
    .b({_al_u4919_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 }),
    .c({_al_u4921_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ,_al_u4920_o}),
    .mi({open_n42941,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .f({_al_u4922_o,_al_u4921_o}),
    .q({open_n42946,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 }));  // ../RTL/cortexm0ds_logic.v(19993)
  EG_PHY_LSLICE #(
    //.LUTF0("(D@(B*~(~C*A)))"),
    //.LUTF1("(A*~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    //.LUTG0("(D@(B*~(~C*A)))"),
    //.LUTG1("(A*~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    .INIT_LUTF0(16'b0011101111000100),
    .INIT_LUTF1(16'b0010000010101000),
    .INIT_LUTG0(16'b0011101111000100),
    .INIT_LUTG1(16'b0010000010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4923|_al_u5615  (
    .a({_al_u4922_o,_al_u4056_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ,_al_u5614_o}),
    .c({_al_u4056_o,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 }),
    .f({_al_u4923_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[16]_i1[16]_o_lutinv }));
  // ../RTL/cortexm0ds_logic.v(19896)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001000111110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4925|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ,open_n42971}),
    .b({_al_u4438_o,open_n42972}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u4925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .q({open_n42989,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 }));  // ../RTL/cortexm0ds_logic.v(19896)
  // ../RTL/cortexm0ds_logic.v(19939)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4926|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ,open_n42990}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ,open_n42991}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhbbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .q({open_n43012,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 }));  // ../RTL/cortexm0ds_logic.v(19939)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(D*~(C@B))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"))
    \_al_u4927|_al_u4933  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 }),
    .f({_al_u4927_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D))"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D))"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000100000101000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000100000101000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4928|_al_u4940  (
    .a({open_n43035,_al_u4927_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }),
    .d({_al_u4927_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 }),
    .f({_al_u4928_o,_al_u4940_o}));
  // ../RTL/cortexm0ds_logic.v(18034)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*A*~(D*~B))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*A*~(D*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b1000000010100000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4929|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6_reg  (
    .a({_al_u4925_o,open_n43060}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ,_al_u5828_o}),
    .c({_al_u4928_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87iu6 ,open_n43079}),
    .q({open_n43083,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 }));  // ../RTL/cortexm0ds_logic.v(18034)
  // ../RTL/cortexm0ds_logic.v(18033)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0100101101001101),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0100101101001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4930|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ,open_n43084}),
    .b({_al_u4438_o,_al_u5826_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .f({_al_u4930_o,open_n43103}),
    .q({open_n43107,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }));  // ../RTL/cortexm0ds_logic.v(18033)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(~D*C*B*~A)"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(~D*C*B*~A)"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b0000000001000000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4932|_al_u4931  (
    .a({_al_u4930_o,open_n43108}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }),
    .c({_al_u4931_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 }),
    .f({_al_u4932_o,_al_u4931_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(A*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1000101000000010),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000101000000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4935|_al_u4974  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 ,_al_u4922_o}),
    .b({_al_u4934_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ,_al_u4056_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 }),
    .f({_al_u4935_o,_al_u4974_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(~D*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~C*~B)*~(~D*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111110001010100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111110001010100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4936|_al_u4941  (
    .a({open_n43157,_al_u4438_o}),
    .b({open_n43158,_al_u4940_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,_al_u4935_o}),
    .d({_al_u4935_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ,_al_u4941_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~B*~(~D*~(~C*~A)))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0011001100000001),
    .MODE("LOGIC"))
    \_al_u4937|_al_u4934  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X87iu6 ,open_n43183}),
    .b({_al_u4932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }),
    .f({_al_u4937_o,_al_u4934_o}));
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4938|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b5  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ,_al_u4121_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u4938_o,\u_cmsdk_mcu/HADDR [7]}),
    .q({open_n43222,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [5]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  // ../RTL/cortexm0ds_logic.v(17859)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("(~D*~C*B*~A)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("(~D*~C*B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4939|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6_reg  (
    .a({_al_u4937_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({_al_u4938_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [5]}),
    .mi({open_n43226,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .f({_al_u4939_o,_al_u5828_o}),
    .q({open_n43242,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 }));  // ../RTL/cortexm0ds_logic.v(17859)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u493|_al_u492  (
    .a({open_n43243,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsubsys_interrupt [1]}),
    .b({_al_u491_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full }),
    .c({_al_u492_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .d({_al_u473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .f({_al_u493_o,_al_u492_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*~(D*B)))"),
    //.LUT1("(~A*~(D*C*~B))"),
    .INIT_LUT0(16'b1010100010100000),
    .INIT_LUT1(16'b0100010101010101),
    .MODE("LOGIC"))
    \_al_u4943|_al_u4942  (
    .a({_al_u4942_o,_al_u4941_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv }),
    .c({_al_u4438_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J17iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 }),
    .f({_al_u4943_o,_al_u4942_o}));
  // ../RTL/cortexm0ds_logic.v(19819)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(D*C*B*~A)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(D*C*B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4944|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6_reg  (
    .a({_al_u4943_o,open_n43288}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ,_al_u5824_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .f({_al_u4944_o,open_n43307}),
    .q({open_n43311,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 }));  // ../RTL/cortexm0ds_logic.v(19819)
  // ../RTL/cortexm0ds_logic.v(18032)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4945|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,_al_u5822_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .f({_al_u4945_o,open_n43332}),
    .q({open_n43336,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 }));  // ../RTL/cortexm0ds_logic.v(18032)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~A*~(~C*~B))"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(D*~A*~(~C*~B))"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b0101010000000000),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0101010000000000),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4946|_al_u4949  (
    .a({open_n43337,_al_u4946_o}),
    .b({_al_u4938_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv }),
    .c({_al_u4945_o,_al_u4438_o}),
    .d({_al_u4438_o,_al_u4948_o}),
    .f({_al_u4946_o,_al_u4949_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B@D))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000110000000011),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4948|_al_u4947  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mz6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 }),
    .c({_al_u4947_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nw6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }),
    .f({_al_u4948_o,_al_u4947_o}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u494|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b0  (
    .b({_al_u493_o,open_n43386}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 }),
    .mi({open_n43390,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u494_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n46 }),
    .q({open_n43405,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [0]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(A*~(D*C*B))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010101010101010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0010101010101010),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4950|u_cmsdk_mcu/u_ahb_ram/reg0_b7  (
    .a({open_n43406,\u_cmsdk_mcu/HADDR [7]}),
    .b({open_n43407,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 }),
    .mi({open_n43411,\u_cmsdk_mcu/HADDR [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4950_o,_al_u6285_o}),
    .q({open_n43426,\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [7]}));  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~A*~(D*~(~C*~B)))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~A*~(D*~(~C*~B)))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000101010101),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4951|_al_u4446  (
    .a({_al_u4939_o,open_n43427}),
    .b({_al_u4944_o,open_n43428}),
    .c({_al_u4949_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 }),
    .d({_al_u4950_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 }),
    .f({_al_u4951_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(D*C*~B*~A)"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0001000000000000),
    .MODE("LOGIC"))
    \_al_u4954|_al_u5817  (
    .a({_al_u4951_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tszhu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv ,_al_u5816_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 ,_al_u4492_o}),
    .d({_al_u4953_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 }),
    .f({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }));
  // ../RTL/cortexm0ds_logic.v(18139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4955|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6_reg  (
    .b({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,_al_u4955_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4955_o,open_n43488}),
    .q({open_n43492,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }));  // ../RTL/cortexm0ds_logic.v(18139)
  // ../RTL/cortexm0ds_logic.v(17977)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4957|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6_reg  (
    .b({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,_al_u4957_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4957_o,open_n43508}),
    .q({open_n43512,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }));  // ../RTL/cortexm0ds_logic.v(17977)
  // ../RTL/cortexm0ds_logic.v(18096)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(A*~(B*~(D@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b0010101010100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4959|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,open_n43513}),
    .b({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ,_al_u4959_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4959_o,open_n43527}),
    .q({open_n43531,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }));  // ../RTL/cortexm0ds_logic.v(18096)
  // ../RTL/cortexm0ds_logic.v(18021)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4961|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,open_n43532}),
    .b({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 ,_al_u4961_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4961_o,open_n43550}),
    .q({open_n43554,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }));  // ../RTL/cortexm0ds_logic.v(18021)
  // ../RTL/cortexm0ds_logic.v(18039)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4963|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,open_n43555}),
    .b({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am6iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,_al_u4963_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4963_o,open_n43569}),
    .q({open_n43573,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }));  // ../RTL/cortexm0ds_logic.v(18039)
  // ../RTL/cortexm0ds_logic.v(18129)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(A*~(B*~(D@C)))"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(A*~(B*~(D@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0010101010100010),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0010101010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4965|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,open_n43574}),
    .b({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({_al_u4438_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ,_al_u4965_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4965_o,open_n43592}),
    .q({open_n43596,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }));  // ../RTL/cortexm0ds_logic.v(18129)
  // ../RTL/cortexm0ds_logic.v(17823)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(A*~(B*~(D@C)))"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(A*~(B*~(D@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0010101010100010),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0010101010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4967|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,open_n43597}),
    .b({_al_u4954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({_al_u4438_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 ,_al_u4967_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u4967_o,open_n43615}),
    .q({open_n43619,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }));  // ../RTL/cortexm0ds_logic.v(17823)
  // ../RTL/cortexm0ds_logic.v(17972)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4969|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6_reg  (
    .a({_al_u4545_o,open_n43620}),
    .b({_al_u4546_o,_al_u3889_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/HADDR[27]_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({_al_u4553_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .mi({open_n43624,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .f({_al_u4969_o,_al_u4553_o}),
    .q({open_n43640,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 }));  // ../RTL/cortexm0ds_logic.v(17972)
  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4970|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b8  (
    .a({_al_u4923_o,open_n43641}),
    .b({_al_u4969_o,_al_u4970_o}),
    .c({\u_cmsdk_mcu/HADDR [12],_al_u4971_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({_al_u4544_o,_al_u4916_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4970_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel }),
    .q({open_n43657,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [8]}));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4971|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b11  (
    .b({\u_cmsdk_mcu/HADDR [14],_al_u4126_o}),
    .c({\u_cmsdk_mcu/HADDR [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4971_o,\u_cmsdk_mcu/HADDR [13]}),
    .q({open_n43679,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [13]}));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4975|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b12  (
    .a({_al_u4973_o,open_n43680}),
    .b({_al_u4974_o,_al_u4131_o}),
    .c({\u_cmsdk_mcu/HADDR [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4975_o,\u_cmsdk_mcu/HADDR [14]}),
    .q({open_n43700,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [14]}));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4977|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b7  (
    .c({_al_u4974_o,_al_u4975_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({_al_u4971_o,_al_u4917_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4977_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/sysctrl_hsel }),
    .q({open_n43720,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [7]}));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~B*~(D*C*A))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0001001100110011),
    .MODE("LOGIC"))
    \_al_u4983|_al_u4982  (
    .a({_al_u695_o,open_n43721}),
    .b({_al_u4982_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }),
    .c({_al_u1582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edapw6_lutinv ,_al_u1266_o}),
    .f({_al_u4983_o,_al_u4982_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~A*~(C*B)))"),
    //.LUTF1("(~D*~C*B*~A)"),
    //.LUTG0("(D*~(~A*~(C*B)))"),
    //.LUTG1("(~D*~C*B*~A)"),
    .INIT_LUTF0(16'b1110101000000000),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b1110101000000000),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4984|_al_u4981  (
    .a({_al_u4981_o,_al_u3618_o}),
    .b({_al_u4983_o,_al_u1346_o}),
    .c({_al_u3187_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 }),
    .d({_al_u3995_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u4984_o,_al_u4981_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~B*~(D*~A)))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b1101000011000000),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u4985|_al_u6817  (
    .a({open_n43766,_al_u3103_o}),
    .b({_al_u2868_o,_al_u1329_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 }),
    .d({_al_u3103_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u4985_o,_al_u6817_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"))
    \_al_u4987|_al_u4986  (
    .a({_al_u3118_o,open_n43787}),
    .b({_al_u4986_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({_al_u1271_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,_al_u1266_o}),
    .f({_al_u4987_o,_al_u4986_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(A*~(~B*~(~D*~C)))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(A*~(~B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b1000100010001010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b1000100010001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4989|_al_u4988  (
    .a({_al_u4984_o,_al_u4985_o}),
    .b({_al_u4988_o,_al_u4987_o}),
    .c({_al_u3103_o,_al_u1269_o}),
    .d({_al_u1342_o,_al_u1342_o}),
    .f({_al_u4989_o,_al_u4988_o}));
  // ../RTL/cortexm0ds_logic.v(18441)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(~D*~B*~A))"),
    //.LUTF1("(C*~(~D*~(B*~A)))"),
    //.LUTG0("~(~C*~(~D*~B*~A))"),
    //.LUTG1("(C*~(~D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110001),
    .INIT_LUTF1(16'b1111000001000000),
    .INIT_LUTG0(16'b1111000011110001),
    .INIT_LUTG1(16'b1111000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4990|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6_reg  (
    .a({_al_u4989_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3xhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u4990_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,_al_u3797_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4990_o,open_n43849}),
    .q({open_n43853,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }));  // ../RTL/cortexm0ds_logic.v(18441)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4992|_al_u4418  (
    .a({open_n43854,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrhiu6 }),
    .b({open_n43855,_al_u3797_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 ,_al_u1809_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z18iu6_lutinv ,_al_u3122_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S18iu6 }));
  // ../RTL/cortexm0ds_logic.v(18054)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u4993|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 ,open_n43876}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 ,_al_u3887_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7cow6 ,_al_u3889_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3436 ),
    .clk(XTAL1_wire),
    .d({_al_u4495_o,_al_u3885_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4993_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7cow6 }),
    .q({open_n43892,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz3qw6 }));  // ../RTL/cortexm0ds_logic.v(18054)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(D*~C*~B*~A)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000000100000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4994|_al_u4546  (
    .a({_al_u3885_o,open_n43893}),
    .b({_al_u3887_o,_al_u3885_o}),
    .c({_al_u3889_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 }),
    .d({_al_u4197_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u4994_o,_al_u4546_o}));
  // ../RTL/cmsdk_mcu_sysctrl.v(250)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u499|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_reg  (
    .a({open_n43918,_al_u497_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe [0],_al_u499_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_write_enable ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_write ),
    .clk(XTAL1_wire),
    .d({_al_u498_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}),
    .mi({open_n43922,\u_cmsdk_mcu/HWDATA [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u499_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_remap_write }),
    .q({open_n43937,\u_cmsdk_mcu/u_cmsdk_mcu_system/remap_ctrl }));  // ../RTL/cmsdk_mcu_sysctrl.v(250)
  // ../RTL/cmsdk_ahb_to_iop.v(105)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(~D*~C*A))"),
    //.LUTF1("(~A*~(~D*C*B))"),
    //.LUTG0("~(B*~(~D*~C*A))"),
    //.LUTG1("(~A*~(~D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100111011),
    .INIT_LUTF1(16'b0101010100010101),
    .INIT_LUTG0(16'b0011001100111011),
    .INIT_LUTG1(16'b0101010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5000|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/IOTRANS_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ,_al_u4993_o}),
    .c({_al_u4994_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7cow6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 ,_al_u4994_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5000_o,\u_cmsdk_mcu/HTRANS [1]}),
    .q({open_n43958,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS }));  // ../RTL/cmsdk_ahb_to_iop.v(105)
  // ../RTL/cmsdk_ahb_to_iop.v(96)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~((D*~C))*~(A)+B*(D*~C)*~(A)+~(B)*(D*~C)*A+B*(D*~C)*A)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100111001000100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5006|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg1_b0  (
    .a({open_n43959,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .b({open_n43960,_al_u4542_o}),
    .c({\u_cmsdk_mcu/HADDR [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzhu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HSIZE [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5006_o,\u_cmsdk_mcu/HSIZE [0]}),
    .q({open_n43977,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [0]}));  // ../RTL/cmsdk_ahb_to_iop.v(96)
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5010|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b0  (
    .c({_al_u5009_o,_al_u5009_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel ,\u_cmsdk_mcu/u_cmsdk_mcu_system/sysctrl_hsel }),
    .mi({open_n43985,\u_cmsdk_mcu/HADDR [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access }),
    .q({open_n44000,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(A*~(~D*~C*~B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(A*~(~D*~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010101010101000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5017|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b4  (
    .a({_al_u4917_o,open_n44001}),
    .b({_al_u4975_o,open_n44002}),
    .c({_al_u4977_o,_al_u4923_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({_al_u4923_o,_al_u4917_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5017_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hsel }),
    .q({open_n44022,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]}));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u5020|_al_u4492  (
    .b({_al_u4492_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5020_o,_al_u4492_o}));
  // ../RTL/cortexm0ds_logic.v(18268)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5021|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6dbx6 }),
    .mi({open_n44048,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .f({_al_u5021_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8liu6 }),
    .q({open_n44064,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 }));  // ../RTL/cortexm0ds_logic.v(18268)
  // ../RTL/cortexm0ds_logic.v(18246)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5023|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,_al_u5730_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,_al_u5759_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dncax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 }),
    .mi({open_n44075,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .f({_al_u5023_o,_al_u5760_o}),
    .q({open_n44080,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krbax6 }));  // ../RTL/cortexm0ds_logic.v(18246)
  // ../RTL/cortexm0ds_logic.v(18290)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5025|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,open_n44081}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv }),
    .mi({open_n44085,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .f({_al_u5025_o,_al_u5782_o}),
    .q({open_n44101,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Widax6 }));  // ../RTL/cortexm0ds_logic.v(18290)
  // ../RTL/cortexm0ds_logic.v(18160)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5026|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6_reg  (
    .a({_al_u5024_o,_al_u2270_o}),
    .b({_al_u5025_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n44112,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .f({_al_u5026_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvow6 }),
    .q({open_n44117,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 }));  // ../RTL/cortexm0ds_logic.v(18160)
  // ../RTL/cortexm0ds_logic.v(17983)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C)*~(A)+~(D*B)*C*~(A)+~(~(D*B))*C*A+~(D*B)*C*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(~(D*B)*~(C)*~(A)+~(D*B)*C*~(A)+~(~(D*B))*C*A+~(D*B)*C*A)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100111000001010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0100111000001010),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5027|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6_reg  (
    .a({open_n44118,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr4iu6_lutinv }),
    .b({open_n44119,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 }),
    .c({_al_u5001_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ur4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,open_n44137}),
    .q({open_n44141,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }));  // ../RTL/cortexm0ds_logic.v(17983)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C*B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(A*~(D*C*B))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b0010101010101010),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0010101010101010),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5028|_al_u5047  (
    .a({open_n44142,_al_u5020_o}),
    .b({_al_u1286_o,_al_u5028_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 }),
    .d({_al_u5026_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .f({_al_u5028_o,_al_u5047_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~A)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(D*~C*~B*~A)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000100000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5030|_al_u540  (
    .a({open_n44167,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .d({_al_u540_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .f({_al_u5030_o,_al_u540_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5032|_al_u5204  (
    .a({_al_u5029_o,open_n44192}),
    .b({_al_u5031_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ,_al_u5031_o}),
    .f({_al_u5032_o,_al_u5204_o}));
  // ../RTL/cortexm0ds_logic.v(19269)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5034|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6_reg  (
    .a({open_n44217,\u_cmsdk_mcu/HWDATA [30]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 }),
    .clk(XTAL1_wire),
    .d({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fllow6_lutinv ,open_n44231}),
    .q({open_n44235,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 }));  // ../RTL/cortexm0ds_logic.v(19269)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~C*~B*D)"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"))
    \_al_u5035|_al_u5033  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5038|_al_u5037  (
    .a({open_n44258,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 }),
    .d({_al_u5037_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 }),
    .f({_al_u5038_o,_al_u5037_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5039|_al_u546  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv }),
    .b({_al_u546_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .f({_al_u5039_o,_al_u546_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5041|_al_u5036  (
    .a({_al_u5036_o,_al_u5032_o}),
    .b({_al_u5038_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fllow6_lutinv }),
    .c({_al_u5039_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .d({_al_u5040_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 ,_al_u5036_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5043|_al_u541  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u540_o}),
    .b({_al_u540_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .c({_al_u1385_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5044|_al_u612  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 }),
    .f({_al_u5044_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5045|_al_u5042  (
    .b({open_n44379,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*~A*~(~D*B))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"))
    \_al_u5049|_al_u5048  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,open_n44404}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 }),
    .c({_al_u5048_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5049_o,_al_u5048_o}));
  // ../RTL/cortexm0ds_logic.v(17963)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5051|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6_reg  (
    .a({_al_u5047_o,open_n44425}),
    .b({_al_u5050_o,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc2qw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 ,_al_u5051_o}),
    .f({_al_u5051_o,open_n44440}),
    .q({open_n44444,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 }));  // ../RTL/cortexm0ds_logic.v(17963)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5052|_al_u5019  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 }),
    .f({_al_u5052_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahwiu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(~C*B)*~(D*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0101000111110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0101000111110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5053|_al_u5308  (
    .a({open_n44471,_al_u5052_o}),
    .b({open_n44472,_al_u5020_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ,_al_u5307_o}),
    .d({_al_u5052_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 }),
    .f({_al_u5053_o,_al_u5308_o}));
  // ../RTL/cortexm0ds_logic.v(18047)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5055|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u5050_o,_al_u1741_o}),
    .f({_al_u5055_o,open_n44513}),
    .q({open_n44517,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 }));  // ../RTL/cortexm0ds_logic.v(18047)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~D*~C*B*A)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"))
    \_al_u5057|_al_u673  (
    .a({_al_u533_o,open_n44518}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ,_al_u533_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv }),
    .f({_al_u5057_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*A*~(D*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*A*~(D*B))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000001000001010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000001000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5058|_al_u5056  (
    .a({_al_u5056_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({_al_u5057_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 }),
    .f({_al_u5058_o,_al_u5056_o}));
  // ../RTL/cortexm0ds_logic.v(17253)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000011110100),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1011000011110100),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5059|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6_reg  (
    .a({open_n44563,_al_u2741_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 }),
    .clk(XTAL1_wire),
    .d({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5059_o,open_n44581}),
    .q({open_n44585,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 }));  // ../RTL/cortexm0ds_logic.v(17253)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5060|_al_u3527  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 }),
    .d({_al_u5059_o,_al_u2741_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 ,_al_u3527_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*~C))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b1000000010001000),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5061|_al_u5062  (
    .a({_al_u5058_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 ,_al_u5061_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u1862_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5061_o,_al_u5062_o}));
  // ../RTL/cortexm0ds_logic.v(18046)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5063|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6_reg  (
    .b({_al_u5020_o,_al_u5053_o}),
    .c({_al_u5062_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 }),
    .clk(XTAL1_wire),
    .d({_al_u5055_o,_al_u5063_o}),
    .f({_al_u5063_o,open_n44648}),
    .q({open_n44652,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rr3qw6 }));  // ../RTL/cortexm0ds_logic.v(18046)
  // ../RTL/cortexm0ds_logic.v(17222)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000011110100),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1011000011110100),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5065|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6_reg  (
    .a({open_n44653,_al_u2733_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 }),
    .clk(XTAL1_wire),
    .d({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwfow6_lutinv ,open_n44671}),
    .q({open_n44675,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usipw6 }));  // ../RTL/cortexm0ds_logic.v(17222)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5066|_al_u3512  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwfow6_lutinv ,_al_u2733_o}),
    .f({_al_u5066_o,_al_u3512_o}));
  // ../RTL/cortexm0ds_logic.v(18407)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D@C))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*A*~(D@C))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000001000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5070|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 ,_al_u5590_o}),
    .b({_al_u5069_o,_al_u5593_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwihu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 }),
    .mi({open_n44705,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .f({_al_u5070_o,_al_u5597_o}),
    .q({open_n44721,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khgax6 }));  // ../RTL/cortexm0ds_logic.v(18407)
  // ../RTL/cortexm0ds_logic.v(18409)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5072|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibqpw6 }),
    .mi({open_n44725,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .f({_al_u5072_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ocniu6 }),
    .q({open_n44741,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 }));  // ../RTL/cortexm0ds_logic.v(18409)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*~(D*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0100000011000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5073|_al_u5071  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({_al_u5071_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({_al_u5072_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 }),
    .f({_al_u5073_o,_al_u5071_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(D*~A))"),
    //.LUT1("(C*A*~(~D*B))"),
    .INIT_LUT0(16'b1000000011000000),
    .INIT_LUT1(16'b1010000000100000),
    .MODE("LOGIC"))
    \_al_u5074|_al_u5320  (
    .a({_al_u5070_o,_al_u4688_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,_al_u5319_o}),
    .c({_al_u5073_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 }),
    .d({_al_u1859_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5074_o,_al_u5320_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5075|_al_u5087  (
    .b({_al_u5074_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ,_al_u5086_o}),
    .d({_al_u5020_o,_al_u5020_o}),
    .f({_al_u5075_o,_al_u5087_o}));
  // ../RTL/cortexm0ds_logic.v(17554)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5076|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqgax6 }),
    .clk(XTAL1_wire),
    .d({_al_u5075_o,_al_u5076_o}),
    .f({_al_u5076_o,open_n44828}),
    .q({open_n44832,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idqpw6 }));  // ../RTL/cortexm0ds_logic.v(17554)
  // ../RTL/cortexm0ds_logic.v(19263)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000011110100),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1011000011110100),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5078|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6_reg  (
    .a({open_n44833,_al_u2729_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 }),
    .clk(XTAL1_wire),
    .d({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5078_o,open_n44851}),
    .q({open_n44855,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 }));  // ../RTL/cortexm0ds_logic.v(19263)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5079|_al_u3507  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 }),
    .d({_al_u5078_o,_al_u2729_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 ,_al_u3507_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u507|_al_u504  (
    .a({open_n44882,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*~(~D*B))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b1010000000100000),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u5080|_al_u5168  (
    .a({open_n44903,_al_u5164_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .c({_al_u1856_o,_al_u5167_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,_al_u1844_o}),
    .f({_al_u5080_o,_al_u5168_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u5082|_al_u5081  (
    .a({open_n44924,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({_al_u5081_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 }),
    .f({_al_u5082_o,_al_u5081_o}));
  // ../RTL/cortexm0ds_logic.v(19965)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5084|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,open_n44945}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,open_n44946}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5084_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .q({open_n44967,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 }));  // ../RTL/cortexm0ds_logic.v(19965)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5085|_al_u5083  (
    .a({open_n44968,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({_al_u5083_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5084_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nybbx6 }),
    .d({_al_u5082_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 }),
    .f({_al_u5085_o,_al_u5083_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5086|_al_u7219  (
    .a({_al_u5080_o,_al_u4289_o}),
    .b({_al_u5085_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [26]}),
    .f({_al_u5086_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zccow6 }));
  // ../RTL/cortexm0ds_logic.v(19942)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5088|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 }),
    .clk(XTAL1_wire),
    .d({_al_u5087_o,_al_u5088_o}),
    .f({_al_u5088_o,open_n45025}),
    .q({open_n45029,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0cbx6 }));  // ../RTL/cortexm0ds_logic.v(19942)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5090|_al_u5171  (
    .b({open_n45032,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 }),
    .d({_al_u5049_o,_al_u5090_o}),
    .f({_al_u5090_o,_al_u5171_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5091|_al_u5310  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 }),
    .d({_al_u5090_o,_al_u5090_o}),
    .f({_al_u5091_o,_al_u5310_o}));
  // ../RTL/cortexm0ds_logic.v(17701)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011000011110100),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5092|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,_al_u2725_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5092_o,open_n45092}),
    .q({open_n45096,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 }));  // ../RTL/cortexm0ds_logic.v(17701)
  // ../RTL/cortexm0ds_logic.v(19949)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5095|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,open_n45097}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n45098}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5095_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .q({open_n45119,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 }));  // ../RTL/cortexm0ds_logic.v(19949)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5099|_al_u5097  (
    .a({open_n45120,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({_al_u5097_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5098_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8cbx6 }),
    .d({_al_u5096_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 }),
    .f({_al_u5099_o,_al_u5097_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5100|_al_u7216  (
    .a({_al_u5094_o,_al_u4289_o}),
    .b({_al_u5099_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [25]}),
    .f({_al_u5100_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhcow6 }));
  // ../RTL/cortexm0ds_logic.v(19954)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(A*~(B*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b1010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5101|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6_reg  (
    .a({_al_u5091_o,open_n45161}),
    .b({_al_u5020_o,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 }),
    .clk(XTAL1_wire),
    .d({_al_u5100_o,_al_u5101_o}),
    .f({_al_u5101_o,open_n45176}),
    .q({open_n45180,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cncbx6 }));  // ../RTL/cortexm0ds_logic.v(19954)
  // ../RTL/cortexm0ds_logic.v(20154)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5103|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6_reg  (
    .b({open_n45183,_al_u5052_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({_al_u5052_o,_al_u5103_o}),
    .mi({open_n45194,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .f({_al_u5103_o,_al_u5104_o}),
    .q({open_n45199,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2ibx6 }));  // ../RTL/cortexm0ds_logic.v(20154)
  // ../RTL/cortexm0ds_logic.v(19257)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011000011110100),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5105|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6_reg  (
    .a({open_n45200,_al_u2721_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 }),
    .clk(XTAL1_wire),
    .d({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5105_o,open_n45214}),
    .q({open_n45218,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 }));  // ../RTL/cortexm0ds_logic.v(19257)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5106|_al_u3497  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 }),
    .d({_al_u5105_o,_al_u2721_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 ,_al_u3497_o}));
  // ../RTL/cortexm0ds_logic.v(18269)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5109|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n45241}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,open_n45242}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .mi({open_n45246,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .f({_al_u5109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 }),
    .q({open_n45262,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 }));  // ../RTL/cortexm0ds_logic.v(18269)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*A)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(D*~C*~B*A)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u510|_al_u512  (
    .a({open_n45263,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }));
  // ../RTL/cortexm0ds_logic.v(17995)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D*~(~C*A)))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~B*~(D*~(~C*A)))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110111001100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111110111001100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5110|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6_reg  (
    .a({_al_u927_o,_al_u927_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u933_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5110_o,open_n45305}),
    .q({open_n45309,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nj2qw6 }));  // ../RTL/cortexm0ds_logic.v(17995)
  // ../RTL/cortexm0ds_logic.v(18179)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5111|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,open_n45310}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n45311}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bp2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5111_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .q({open_n45328,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 }));  // ../RTL/cortexm0ds_logic.v(18179)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5112|_al_u5108  (
    .a({_al_u5108_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u5109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .c({_al_u5110_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 }),
    .d({_al_u5111_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 }),
    .f({_al_u5112_o,_al_u5108_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5113|_al_u7213  (
    .a({_al_u5107_o,_al_u4289_o}),
    .b({_al_u5112_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [24]}),
    .f({_al_u5113_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmcow6 }));
  // ../RTL/cortexm0ds_logic.v(17997)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*A*~(D*C))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110111011101),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5114|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6_reg  (
    .a({open_n45377,_al_u5104_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ,_al_u5114_o}),
    .c({_al_u5113_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5020_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 }),
    .f({_al_u5114_o,open_n45392}),
    .q({open_n45396,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fl2qw6 }));  // ../RTL/cortexm0ds_logic.v(17997)
  // ../RTL/cortexm0ds_logic.v(18270)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5116|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n45397}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,open_n45398}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5116_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .q({open_n45419,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 }));  // ../RTL/cortexm0ds_logic.v(18270)
  // ../RTL/cortexm0ds_logic.v(18314)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A*(C@B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010000000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5117|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6_reg  (
    .a({open_n45420,_al_u5787_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u4184_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5116_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 }),
    .mi({open_n45431,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .f({_al_u5117_o,_al_u5788_o}),
    .q({open_n45436,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jieax6 }));  // ../RTL/cortexm0ds_logic.v(18314)
  // ../RTL/cortexm0ds_logic.v(18180)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5118|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6_reg  (
    .a({_al_u927_o,open_n45437}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrihu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uh2qw6 ,_al_u5599_o}),
    .mi({open_n45441,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .f({_al_u5118_o,_al_u5603_o}),
    .q({open_n45457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6aax6 }));  // ../RTL/cortexm0ds_logic.v(18180)
  // ../RTL/cortexm0ds_logic.v(20159)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101110001010),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1011101110001010),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5119|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6_reg  (
    .a({open_n45458,_al_u5515_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ,_al_u5516_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5118_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5119_o,open_n45476}),
    .q({open_n45480,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4ibx6 }));  // ../RTL/cortexm0ds_logic.v(20159)
  // ../RTL/cortexm0ds_logic.v(18349)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5121|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ,open_n45481}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgkbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .mi({open_n45492,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5121_o,_al_u5519_o}),
    .q({open_n45496,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 }));  // ../RTL/cortexm0ds_logic.v(18349)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5122|_al_u5120  (
    .a({_al_u5117_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u5119_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({_al_u5120_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 }),
    .d({_al_u5121_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 }),
    .f({_al_u5122_o,_al_u5120_o}));
  // ../RTL/cortexm0ds_logic.v(17316)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~C*~(D)*~((B*~A))+~C*D*~((B*~A))+~(~C)*D*(B*~A)+~C*D*(B*~A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000011110100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1011000011110100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5123|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,_al_u2717_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgeow6 ,open_n45538}),
    .q({open_n45542,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 }));  // ../RTL/cortexm0ds_logic.v(17316)
  // ../RTL/cortexm0ds_logic.v(17307)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110001010),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5125|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ,_al_u5637_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u5638_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5125_o,open_n45556}),
    .q({open_n45560,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpkpw6 }));  // ../RTL/cortexm0ds_logic.v(17307)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*C*B))"),
    //.LUT1("(C*B*~(~D*A))"),
    .INIT_LUT0(16'b0010101010101010),
    .INIT_LUT1(16'b1100000001000000),
    .MODE("LOGIC"))
    \_al_u5126|_al_u5127  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,_al_u5020_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .c({_al_u5125_o,_al_u5122_o}),
    .d({_al_u1850_o,_al_u5126_o}),
    .f({_al_u5126_o,_al_u5127_o}));
  // ../RTL/cortexm0ds_logic.v(17309)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*A*~(D*C))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(~B*A*~(D*C))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110111011101),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1111110111011101),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5128|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6_reg  (
    .a({open_n45581,_al_u5128_o}),
    .b({_al_u5052_o,_al_u5103_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/No3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5127_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 }),
    .f({_al_u5128_o,open_n45600}),
    .q({open_n45604,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrkpw6 }));  // ../RTL/cortexm0ds_logic.v(17309)
  // ../RTL/cortexm0ds_logic.v(20018)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5130|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tlebx6 }),
    .mi({open_n45615,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .f({_al_u5130_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ctliu6 }),
    .q({open_n45620,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 }));  // ../RTL/cortexm0ds_logic.v(20018)
  // ../RTL/cortexm0ds_logic.v(20017)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5131|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6_reg  (
    .a({open_n45621,_al_u1952_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5130_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n45632,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .f({_al_u5131_o,_al_u2237_o}),
    .q({open_n45637,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 }));  // ../RTL/cortexm0ds_logic.v(20017)
  // ../RTL/cortexm0ds_logic.v(20016)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*(D@C))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(B*A*(D@C))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000100010000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5133|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u5806_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,_al_u5807_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 ,_al_u4086_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 }),
    .mi({open_n45641,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .f({_al_u5133_o,_al_u5808_o}),
    .q({open_n45657,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kpfbx6 }));  // ../RTL/cortexm0ds_logic.v(20016)
  // ../RTL/cortexm0ds_logic.v(20013)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5134|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,open_n45658}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n45659}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5134_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .q({open_n45680,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 }));  // ../RTL/cortexm0ds_logic.v(20013)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(~C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(~C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0011000111110101),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0011000111110101),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5135|_al_u5132  (
    .a({_al_u5131_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .b({_al_u5132_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .c({_al_u5133_o,_al_u1846_o}),
    .d({_al_u5134_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] }),
    .f({_al_u5135_o,_al_u5132_o}));
  // ../RTL/cortexm0ds_logic.v(20037)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5136|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [22]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5136_o,open_n45718}),
    .q({open_n45722,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3gbx6 }));  // ../RTL/cortexm0ds_logic.v(20037)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5137|_al_u1304  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ,open_n45723}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .f({_al_u5137_o,_al_u1304_o}));
  // ../RTL/cortexm0ds_logic.v(20069)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5138|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6_reg  (
    .a({_al_u5136_o,open_n45748}),
    .b({_al_u5137_o,\u_cmsdk_mcu/sram_hrdata [22]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ,\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ,\u_cmsdk_mcu/HWDATA [22]}),
    .mi({open_n45759,\u_cmsdk_mcu/HWDATA [22]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5138_o,\u_cmsdk_mcu/u_ahb_ram/n13 [22]}),
    .q({open_n45763,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 }));  // ../RTL/cortexm0ds_logic.v(20069)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000001110111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5139|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b13  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ,\u_cmsdk_mcu/HWDATA [13]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 }),
    .mi({open_n45774,\u_cmsdk_mcu/HWDATA [13]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5139_o,_al_u3348_o}),
    .q({open_n45778,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [13]}));  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5140|_al_u5261  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ,open_n45779}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 ,_al_u5260_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .f({_al_u5140_o,_al_u5261_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u5142|_al_u3465  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ,open_n45804}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V73bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ,\u_cmsdk_mcu/HWDATA [19]}),
    .f({_al_u5142_o,_al_u3465_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5143|_al_u5141  (
    .a({_al_u5139_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 }),
    .b({_al_u5140_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 }),
    .c({_al_u5141_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 }),
    .d({_al_u5142_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 }),
    .f({_al_u5143_o,_al_u5141_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5144|_al_u3470  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ,open_n45845}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ,\u_cmsdk_mcu/HWDATA [20]}),
    .f({_al_u5144_o,_al_u3470_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u5145|_al_u3448  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ,open_n45870}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ,\u_cmsdk_mcu/HWDATA [17]}),
    .f({_al_u5145_o,_al_u3448_o}));
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000001110111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0010000001110111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5147|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b11  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ,\u_cmsdk_mcu/HWDATA [11]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 }),
    .mi({open_n45894,\u_cmsdk_mcu/HWDATA [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5147_o,_al_u3345_o}),
    .q({open_n45909,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [11]}));  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5148|_al_u5146  (
    .a({_al_u5144_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 }),
    .b({_al_u5145_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 }),
    .c({_al_u5146_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 }),
    .d({_al_u5147_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 }),
    .f({_al_u5148_o,_al_u5146_o}));
  // ../RTL/cortexm0ds_logic.v(20045)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5150|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,open_n45930}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ,open_n45931}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .mi({open_n45935,\u_cmsdk_mcu/HWDATA [22]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zpkow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 }),
    .q({open_n45951,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D7gbx6 }));  // ../RTL/cortexm0ds_logic.v(20045)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5152|_al_u5151  (
    .a({open_n45952,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zpkow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 }),
    .c({_al_u5151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 }),
    .d({_al_u5149_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 }),
    .f({_al_u5152_o,_al_u5151_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*C*B))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0010101010101010),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5155|_al_u5156  (
    .a({_al_u5138_o,_al_u5020_o}),
    .b({_al_u5152_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .c({_al_u5153_o,_al_u5135_o}),
    .d({_al_u5154_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 ,_al_u5156_o}));
  // ../RTL/cortexm0ds_logic.v(20020)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5157|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6_reg  (
    .a({_al_u5156_o,open_n45997}),
    .b({_al_u5090_o,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 ,_al_u5157_o}),
    .f({_al_u5157_o,open_n46016}),
    .q({open_n46020,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 }));  // ../RTL/cortexm0ds_logic.v(20020)
  // ../RTL/cortexm0ds_logic.v(19973)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5159|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u5090_o,_al_u1716_o}),
    .f({_al_u5159_o,open_n46041}),
    .q({open_n46045,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sddbx6 }));  // ../RTL/cortexm0ds_logic.v(19973)
  // ../RTL/cortexm0ds_logic.v(19245)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5160|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [21]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdfow6 ,open_n46059}),
    .q({open_n46063,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 }));  // ../RTL/cortexm0ds_logic.v(19245)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5161|_al_u5227  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdfow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9mow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fdfow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9mow6 }));
  // ../RTL/cortexm0ds_logic.v(17299)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5162|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,_al_u2235_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fdfow6 ,_al_u2228_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 ,\u_cmsdk_mcu/HWDATA [21]}),
    .q({open_n46108,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhkpw6 }));  // ../RTL/cortexm0ds_logic.v(17299)
  // ../RTL/cortexm0ds_logic.v(19992)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5163|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n46109}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n46110}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5163_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .q({open_n46131,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 }));  // ../RTL/cortexm0ds_logic.v(19992)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5164|_al_u5200  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u5163_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 }),
    .f({_al_u5164_o,_al_u5200_o}));
  // ../RTL/cortexm0ds_logic.v(19988)
  EG_PHY_MSLICE #(
    //.LUT0("(C@D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111110000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5165|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,open_n46156}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,open_n46157}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2ebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snihu6 }),
    .mi({open_n46168,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .f({_al_u5165_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[21]_i1[21]_o_lutinv }),
    .q({open_n46173,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6ebx6 }));  // ../RTL/cortexm0ds_logic.v(19988)
  // ../RTL/cortexm0ds_logic.v(19989)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*~A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*C)*~(B*~A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101110111011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000101110111011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5166|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u1943_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n46177,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .f({_al_u5166_o,_al_u2228_o}),
    .q({open_n46193,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 }));  // ../RTL/cortexm0ds_logic.v(19989)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*A*~(D*B))"),
    //.LUTF1("(C*B*~(D*A))"),
    //.LUTG0("(C*A*~(D*B))"),
    //.LUTG1("(C*B*~(D*A))"),
    .INIT_LUTF0(16'b0010000010100000),
    .INIT_LUTF1(16'b0100000011000000),
    .INIT_LUTG0(16'b0010000010100000),
    .INIT_LUTG1(16'b0100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5167|_al_u5024  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u5021_o}),
    .b({_al_u5165_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .c({_al_u5166_o,_al_u5023_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] }),
    .f({_al_u5167_o,_al_u5024_o}));
  // ../RTL/cortexm0ds_logic.v(19994)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(A*~(B*~(D*C)))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(A*~(B*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b1010001000100010),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b1010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5169|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6_reg  (
    .a({_al_u5159_o,open_n46218}),
    .b({_al_u5020_o,_al_u5053_o}),
    .c({_al_u5168_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ,_al_u5169_o}),
    .f({_al_u5169_o,open_n46237}),
    .q({open_n46241,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jhebx6 }));  // ../RTL/cortexm0ds_logic.v(19994)
  // ../RTL/cortexm0ds_logic.v(19239)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5172|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [20]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fe2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrfow6 ,open_n46255}),
    .q({open_n46259,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mp0bx6 }));  // ../RTL/cortexm0ds_logic.v(19239)
  // ../RTL/cortexm0ds_logic.v(17230)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5173|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,_al_u1934_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mrfow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qoyow6 }),
    .f({_al_u5173_o,\u_cmsdk_mcu/HWDATA [20]}),
    .q({open_n46278,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6jpw6 }));  // ../RTL/cortexm0ds_logic.v(17230)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5174|_al_u5176  (
    .a({open_n46279,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcuiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .d({_al_u5173_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 ,_al_u5176_o}));
  // ../RTL/cortexm0ds_logic.v(19981)
  EG_PHY_MSLICE #(
    //.LUT0("((C@B)*(D@A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010000101000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5178|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,_al_u4076_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,_al_u4141_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 }),
    .mi({open_n46310,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .f({_al_u5178_o,_al_u5779_o}),
    .q({open_n46315,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsdbx6 }));  // ../RTL/cortexm0ds_logic.v(19981)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u517|_al_u516  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 ,_al_u374_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(~C*A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0011000111110101),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5180|_al_u5177  (
    .a({_al_u5176_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .b({_al_u5177_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .c({_al_u5178_o,_al_u1841_o}),
    .d({_al_u5179_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] }),
    .f({_al_u5180_o,_al_u5177_o}));
  // ../RTL/cortexm0ds_logic.v(19984)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(A*~(B*~(D*C)))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(A*~(B*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b1010001000100010),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b1010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5181|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6_reg  (
    .a({_al_u5171_o,open_n46358}),
    .b({_al_u5020_o,_al_u5053_o}),
    .c({_al_u5180_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ,_al_u5181_o}),
    .f({_al_u5181_o,open_n46377}),
    .q({open_n46381,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 }));  // ../RTL/cortexm0ds_logic.v(19984)
  // ../RTL/cortexm0ds_logic.v(19233)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5183|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [19]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5183_o,open_n46395}),
    .q({open_n46399,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 }));  // ../RTL/cortexm0ds_logic.v(19233)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5185|_al_u5184  (
    .a({open_n46400,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({_al_u5183_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5jow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 }),
    .d({_al_u5031_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5jow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5187|_al_u5186  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({_al_u5186_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 }),
    .f({_al_u5187_o,_al_u5186_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5190|_al_u7077  (
    .a({open_n46441,_al_u4289_o}),
    .b({_al_u1385_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [18]}),
    .f({_al_u5190_o,_al_u7077_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5191|_al_u5189  (
    .a({_al_u5187_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u5188_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5189_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 }),
    .d({_al_u5190_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6kbx6 }),
    .f({_al_u5191_o,_al_u5189_o}));
  // ../RTL/cortexm0ds_logic.v(20210)
  EG_PHY_MSLICE #(
    //.LUT0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUT1("(D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100000001),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5192|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6_reg  (
    .a({open_n46490,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({_al_u1839_o,_al_u1839_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5191_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 }),
    .f({_al_u5192_o,open_n46505}),
    .q({open_n46509,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vqjbx6 }));  // ../RTL/cortexm0ds_logic.v(20210)
  // ../RTL/cortexm0ds_logic.v(17773)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5194|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6_reg  (
    .a({_al_u5193_o,open_n46510}),
    .b({_al_u5050_o,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 ,_al_u5194_o}),
    .f({_al_u5194_o,open_n46529}),
    .q({open_n46533,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 }));  // ../RTL/cortexm0ds_logic.v(17773)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5197|_al_u5196  (
    .a({open_n46534,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 }),
    .d({_al_u5196_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 }),
    .f({_al_u5197_o,_al_u5196_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*~B*A)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"))
    \_al_u5201|_al_u5199  (
    .a({_al_u5197_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({_al_u5198_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5199_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 }),
    .d({_al_u5200_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Syjbx6 }),
    .f({_al_u5201_o,_al_u5199_o}));
  // ../RTL/cortexm0ds_logic.v(19227)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5202|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6_reg  (
    .a({open_n46579,\u_cmsdk_mcu/HWDATA [18]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 }),
    .clk(XTAL1_wire),
    .d({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbpow6_lutinv ,open_n46593}),
    .q({open_n46597,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 }));  // ../RTL/cortexm0ds_logic.v(19227)
  // ../RTL/cortexm0ds_logic.v(17828)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5205|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6_reg  (
    .a({_al_u5203_o,open_n46598}),
    .b({_al_u5204_o,_al_u2208_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 ,_al_u2201_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 ,\u_cmsdk_mcu/HWDATA [18]}),
    .q({open_n46615,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lywpw6 }));  // ../RTL/cortexm0ds_logic.v(17828)
  // ../RTL/cortexm0ds_logic.v(20211)
  EG_PHY_MSLICE #(
    //.LUT0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUT1("(B*A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100000001),
    .INIT_LUT1(16'b1000000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5206|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6_reg  (
    .a({_al_u5201_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 ,_al_u1836_o}),
    .c({_al_u1836_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 }),
    .f({_al_u5206_o,open_n46630}),
    .q({open_n46634,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usjbx6 }));  // ../RTL/cortexm0ds_logic.v(20211)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*~(D*~B)))"),
    //.LUT1("(A*~(C*~(D*~B)))"),
    .INIT_LUT0(16'b0010101000001010),
    .INIT_LUT1(16'b0010101000001010),
    .MODE("LOGIC"))
    \_al_u5207|_al_u5193  (
    .a({_al_u5020_o,_al_u5020_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa5iu6 ,_al_u4284_o}),
    .c({_al_u5206_o,_al_u5192_o}),
    .d({_al_u927_o,_al_u927_o}),
    .f({_al_u5207_o,_al_u5193_o}));
  // ../RTL/cortexm0ds_logic.v(17825)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5208|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6_reg  (
    .a({_al_u5207_o,open_n46655}),
    .b({_al_u5049_o,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl3qw6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 ,_al_u5208_o}),
    .f({_al_u5208_o,open_n46670}),
    .q({open_n46674,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 }));  // ../RTL/cortexm0ds_logic.v(17825)
  // ../RTL/cortexm0ds_logic.v(19185)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5210|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [11]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fviow6 ,open_n46688}),
    .q({open_n46692,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 }));  // ../RTL/cortexm0ds_logic.v(19185)
  // ../RTL/cortexm0ds_logic.v(17422)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~A*~(~C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110101110),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5212|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6_reg  (
    .a({open_n46693,_al_u2055_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,_al_u1892_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 ,_al_u2062_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yuiow6 ,_al_u2063_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 ,\u_cmsdk_mcu/HWDATA [11]}),
    .q({open_n46710,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofmpw6 }));  // ../RTL/cortexm0ds_logic.v(17422)
  // ../RTL/cortexm0ds_logic.v(19807)
  EG_PHY_LSLICE #(
    //.LUTF0("((C@B)*(D@A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("((C@B)*(D@A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010000101000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010000101000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5213|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,_al_u4116_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u4197_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 }),
    .mi({open_n46714,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .f({_al_u5213_o,_al_u5807_o}),
    .q({open_n46730,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N19bx6 }));  // ../RTL/cortexm0ds_logic.v(19807)
  // ../RTL/cortexm0ds_logic.v(19805)
  EG_PHY_MSLICE #(
    //.LUT0("~(D@(B*~(~C*A)))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010000111011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5214|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 ,_al_u4116_o}),
    .b({_al_u5213_o,_al_u5592_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,_al_u5523_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 }),
    .mi({open_n46741,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .f({_al_u5214_o,_al_u5593_o}),
    .q({open_n46746,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ux8bx6 }));  // ../RTL/cortexm0ds_logic.v(19805)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5215|_al_u7180  (
    .a({open_n46747,_al_u4289_o}),
    .b({_al_u1385_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [10]}),
    .f({_al_u5215_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eriow6 }));
  // ../RTL/cortexm0ds_logic.v(19808)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5216|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,open_n46772}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,open_n46773}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C07bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .mi({open_n46777,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .f({_al_u5216_o,_al_u2063_o}),
    .q({open_n46793,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 }));  // ../RTL/cortexm0ds_logic.v(19808)
  // ../RTL/cortexm0ds_logic.v(19804)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5217|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,open_n46794}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n46795}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5217_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .q({open_n46812,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 }));  // ../RTL/cortexm0ds_logic.v(19804)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(C*~(D*~B)))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(A*~(C*~(D*~B)))"),
    //.LUTG1("(D*C*~B*A)"),
    .INIT_LUTF0(16'b0010101000001010),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0010101000001010),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5218|_al_u5219  (
    .a({_al_u5214_o,_al_u5020_o}),
    .b({_al_u5215_o,_al_u4796_o}),
    .c({_al_u5216_o,_al_u5218_o}),
    .d({_al_u5217_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5218_o,_al_u5219_o}));
  // ../RTL/cortexm0ds_logic.v(19762)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5220|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 }),
    .clk(XTAL1_wire),
    .d({_al_u5219_o,_al_u5220_o}),
    .f({_al_u5220_o,open_n46857}),
    .q({open_n46861,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 }));  // ../RTL/cortexm0ds_logic.v(19762)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u5222|_al_u7174  (
    .a({open_n46862,_al_u4289_o}),
    .b({_al_u1385_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [9]}),
    .f({_al_u5222_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0mow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*~D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"))
    \_al_u5225|_al_u5224  (
    .a({open_n46883,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .b({_al_u5223_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 }),
    .c({_al_u5224_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 }),
    .d({_al_u5222_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 }),
    .f({_al_u5225_o,_al_u5224_o}));
  // ../RTL/cortexm0ds_logic.v(19179)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000011111000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111000011111000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5226|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [10]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9mow6 ,open_n46921}),
    .q({open_n46925,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 }));  // ../RTL/cortexm0ds_logic.v(19179)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5228|_al_u5690  (
    .a({open_n46926,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tptpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9mow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wnxax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ,_al_u5690_o}));
  // ../RTL/cortexm0ds_logic.v(18277)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5229|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwxpw6 }),
    .mi({open_n46950,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .f({_al_u5229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ivmiu6 }),
    .q({open_n46966,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 }));  // ../RTL/cortexm0ds_logic.v(18277)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u522|_al_u5067  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5eiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ,_al_u5067_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5231|_al_u5230  (
    .a({_al_u5225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({_al_u5229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 }),
    .d({_al_u5230_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 }),
    .f({_al_u5231_o,_al_u5230_o}));
  // ../RTL/cortexm0ds_logic.v(17856)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5233|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4ypw6 }),
    .clk(XTAL1_wire),
    .d({_al_u5232_o,_al_u5233_o}),
    .f({_al_u5233_o,open_n47031}),
    .q({open_n47035,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 }));  // ../RTL/cortexm0ds_logic.v(17856)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5235|_al_u7177  (
    .a({open_n47036,_al_u4289_o}),
    .b({_al_u1385_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [8]}),
    .f({_al_u5235_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdjow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5236|_al_u5188  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 }),
    .f({_al_u5236_o,_al_u5188_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*~D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"))
    \_al_u5238|_al_u5237  (
    .a({open_n47085,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .b({_al_u5236_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5237_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 }),
    .d({_al_u5235_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kn1qw6 }),
    .f({_al_u5238_o,_al_u5237_o}));
  // ../RTL/cortexm0ds_logic.v(20206)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000011111000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0111000011111000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5241|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [9]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5241_o,open_n47123}),
    .q({open_n47127,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 }));  // ../RTL/cortexm0ds_logic.v(20206)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5242|_al_u5244  (
    .a({open_n47128,_al_u5242_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ,_al_u5243_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .d({_al_u5241_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 }),
    .f({_al_u5242_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 }));
  // ../RTL/cortexm0ds_logic.v(20208)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~A*~(~C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110101110),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5243|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6_reg  (
    .a({open_n47149,_al_u1971_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,_al_u1892_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5031_o,_al_u1979_o}),
    .f({_al_u5243_o,\u_cmsdk_mcu/HWDATA [9]}),
    .q({open_n47166,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmjbx6 }));  // ../RTL/cortexm0ds_logic.v(20208)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(C*B*~(D*~A))"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b1000000011000000),
    .MODE("LOGIC"))
    \_al_u5245|_al_u6871  (
    .a({_al_u4756_o,_al_u4756_o}),
    .b({_al_u5240_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibsiu6 ,_al_u6819_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u5245_o,_al_u6871_o}));
  // ../RTL/cortexm0ds_logic.v(17942)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("(~(D*B)*~(~C*A))"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b0011000111110101),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b0011000111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5246|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6_reg  (
    .a({_al_u5020_o,open_n47187}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u1687_o}),
    .c({_al_u5245_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .f({_al_u5246_o,open_n47206}),
    .q({open_n47210,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 }));  // ../RTL/cortexm0ds_logic.v(17942)
  // ../RTL/cortexm0ds_logic.v(19173)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5248|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [8]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzdow6 ,open_n47224}),
    .q({open_n47228,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 }));  // ../RTL/cortexm0ds_logic.v(19173)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5250|_al_u5249  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rq0qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wydow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzdow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wydow6 }));
  // ../RTL/cortexm0ds_logic.v(18278)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5251|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n47251}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,open_n47252}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gc1qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5251_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .q({open_n47273,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5dax6 }));  // ../RTL/cortexm0ds_logic.v(18278)
  // ../RTL/cortexm0ds_logic.v(18188)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5252|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 ,open_n47274}),
    .b({_al_u5251_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6ihu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 ,_al_u5539_o}),
    .mi({open_n47278,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .f({_al_u5252_o,_al_u5544_o}),
    .q({open_n47294,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlaax6 }));  // ../RTL/cortexm0ds_logic.v(18188)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u5253|_al_u7183  (
    .a({open_n47295,_al_u4289_o}),
    .b({_al_u1385_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [7]}),
    .f({_al_u5253_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvdow6 }));
  // ../RTL/cortexm0ds_logic.v(18300)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*(D@C))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(B*A*(D@C))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000100010000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5254|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,_al_u5766_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u5767_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N61qw6 ,_al_u4106_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 }),
    .mi({open_n47319,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .f({_al_u5254_o,_al_u5768_o}),
    .q({open_n47335,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1eax6 }));  // ../RTL/cortexm0ds_logic.v(18300)
  // ../RTL/cortexm0ds_logic.v(18170)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5255|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,open_n47336}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n47337}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .mi({open_n47341,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .f({_al_u5255_o,_al_u1902_o}),
    .q({open_n47357,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 }));  // ../RTL/cortexm0ds_logic.v(18170)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*~(D*~B)))"),
    //.LUT1("(D*C*~B*A)"),
    .INIT_LUT0(16'b0010101000001010),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"))
    \_al_u5256|_al_u5257  (
    .a({_al_u5252_o,_al_u5020_o}),
    .b({_al_u5253_o,_al_u4836_o}),
    .c({_al_u5254_o,_al_u5256_o}),
    .d({_al_u5255_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5256_o,_al_u5257_o}));
  // ../RTL/cortexm0ds_logic.v(17937)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5258|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u1685_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u5257_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .f({_al_u5258_o,open_n47394}),
    .q({open_n47398,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qa1qw6 }));  // ../RTL/cortexm0ds_logic.v(17937)
  // ../RTL/cortexm0ds_logic.v(19647)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5262|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ,open_n47399}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ,open_n47400}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ,_al_u2480_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n47404,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5262_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n158 }),
    .q({open_n47419,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 }));  // ../RTL/cortexm0ds_logic.v(19647)
  // ../RTL/cortexm0ds_logic.v(19167)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5263|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6_reg  (
    .a({_al_u5261_o,\u_cmsdk_mcu/HWDATA [7]}),
    .b({_al_u5262_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5263_o,open_n47433}),
    .q({open_n47437,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 }));  // ../RTL/cortexm0ds_logic.v(19167)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5266|_al_u5264  (
    .a({open_n47438,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({_al_u5264_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 }),
    .c({_al_u5265_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 }),
    .d({_al_u5263_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thxax6 }),
    .f({_al_u5266_o,_al_u5264_o}));
  // ../RTL/cortexm0ds_logic.v(19683)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5267|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ,open_n47459}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,open_n47460}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }),
    .mi({open_n47471,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5267_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 }),
    .q({open_n47475,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 }));  // ../RTL/cortexm0ds_logic.v(19683)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5269|_al_u5268  (
    .a({open_n47476,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 }),
    .b({_al_u5267_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .c({_al_u5268_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 }),
    .d({_al_u5266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 ,_al_u5268_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5271|_al_u5270  (
    .a({open_n47501,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .f({_al_u5271_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5273|_al_u611  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ,open_n47528}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqriu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~D*~(~A*~(C*B)))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~D*~(~A*~(C*B)))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011101010),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5274|_al_u374  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqriu6 ,open_n47553}),
    .b({_al_u374_o,open_n47554}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .f({_al_u5274_o,_al_u374_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~(~A*~(D*B)))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1110000010100000),
    .MODE("LOGIC"))
    \_al_u5276|_al_u5275  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ,open_n47579}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ,open_n47580}),
    .c({_al_u5275_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .f({_al_u5276_o,_al_u5275_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*A))"),
    //.LUT1("(~C*~B*D)"),
    .INIT_LUT0(16'b0101111100010011),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"))
    \_al_u5277|_al_u5272  (
    .a({open_n47601,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .b({_al_u5274_o,_al_u5271_o}),
    .c({_al_u5276_o,_al_u1385_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 }));
  // ../RTL/cortexm0ds_logic.v(18279)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5278|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n47622}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,open_n47623}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1mpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5278_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 }),
    .q({open_n47644,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 }));  // ../RTL/cortexm0ds_logic.v(18279)
  // ../RTL/cortexm0ds_logic.v(18091)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u527|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6_reg  (
    .a({_al_u526_o,open_n47645}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 }),
    .mi({open_n47649,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .q({open_n47665,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 }));  // ../RTL/cortexm0ds_logic.v(18091)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~A*~(~D*C*B))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~A*~(~D*C*B))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0101010100010101),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0101010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5281|_al_u5280  (
    .a({_al_u5280_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ,_al_u5280_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*B))"),
    //.LUT1("(C*A*~(D*B))"),
    .INIT_LUT0(16'b0001000001010000),
    .INIT_LUT1(16'b0010000010100000),
    .MODE("LOGIC"))
    \_al_u5282|_al_u5296  (
    .a({_al_u5278_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ,_al_u5295_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk9bx6 }),
    .f({_al_u5282_o,_al_u5296_o}));
  // ../RTL/cortexm0ds_logic.v(18189)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(D@B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*~A*~(D@B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5284|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,_al_u5556_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5ihu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 ,_al_u5519_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 }),
    .mi({open_n47713,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 }),
    .f({_al_u5284_o,_al_u5558_o}),
    .q({open_n47729,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnaax6 }));  // ../RTL/cortexm0ds_logic.v(18189)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(C*B*~(D*A))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0100000011000000),
    .MODE("LOGIC"))
    \_al_u5285|_al_u7200  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsriu6 ,_al_u4290_o}),
    .c({_al_u5284_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [6]}),
    .f({_al_u5285_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W48ow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(C*~(D*~B)))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(A*~(C*~(D*~B)))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0010101000001010),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0010101000001010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5286|_al_u5287  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 ,_al_u5020_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ,_al_u4735_o}),
    .c({_al_u5282_o,_al_u5286_o}),
    .d({_al_u5285_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5286_o,_al_u5287_o}));
  // ../RTL/cortexm0ds_logic.v(20246)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5288|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 }),
    .clk(XTAL1_wire),
    .d({_al_u5287_o,_al_u5288_o}),
    .f({_al_u5288_o,open_n47794}),
    .q({open_n47798,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nckbx6 }));  // ../RTL/cortexm0ds_logic.v(20246)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5292|_al_u535  (
    .c({_al_u5291_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lariu6 ,_al_u533_o}),
    .f({_al_u5292_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u5293|_al_u7197  (
    .a({_al_u5292_o,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u4290_o}),
    .c({_al_u1385_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [5]}),
    .f({_al_u5293_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkeow6 }));
  // ../RTL/cortexm0ds_logic.v(19818)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5294|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n47843}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n47844}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5294_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 }),
    .q({open_n47861,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl9bx6 }));  // ../RTL/cortexm0ds_logic.v(19818)
  // ../RTL/cortexm0ds_logic.v(19816)
  EG_PHY_MSLICE #(
    //.LUT0("((D@B)*(C@A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001001001000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5295|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u4066_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4141_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmeax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 }),
    .mi({open_n47872,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 }),
    .f({_al_u5295_o,_al_u5803_o}),
    .q({open_n47877,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hi9bx6 }));  // ../RTL/cortexm0ds_logic.v(19816)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5298|_al_u5297  (
    .a({_al_u5293_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({_al_u5294_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .c({_al_u5296_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 }),
    .d({_al_u5297_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 }),
    .f({_al_u5298_o,_al_u5297_o}));
  // ../RTL/cortexm0ds_logic.v(19844)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5299|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,open_n47898}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ,open_n47899}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 ,_al_u2478_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n47910,\u_cmsdk_mcu/HWDATA [6]}),
    .f({_al_u5299_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n201 }),
    .q({open_n47915,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ox9bx6 }));  // ../RTL/cortexm0ds_logic.v(19844)
  // ../RTL/cortexm0ds_logic.v(19836)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5301|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [6]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5301_o,open_n47929}),
    .q({open_n47933,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 }));  // ../RTL/cortexm0ds_logic.v(19836)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5303|_al_u5302  (
    .a({_al_u5301_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 }),
    .b({_al_u5302_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 }),
    .f({_al_u5303_o,_al_u5302_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5306|_al_u5304  (
    .a({_al_u5300_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }),
    .b({_al_u5303_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({_al_u5304_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 }),
    .d({_al_u5305_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 ,_al_u5304_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(C*B*~(D*~A))"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b1000000011000000),
    .MODE("LOGIC"))
    \_al_u5307|_al_u6950  (
    .a({_al_u4712_o,_al_u4712_o}),
    .b({_al_u5298_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkriu6 ,_al_u6819_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u5307_o,_al_u6950_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5311|_al_u7159  (
    .a({open_n48002,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] }),
    .d({_al_u5292_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [4]}),
    .f({_al_u5311_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xneow6 }));
  // ../RTL/cortexm0ds_logic.v(19161)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5312|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [5]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5312_o,open_n48036}),
    .q({open_n48040,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 }));  // ../RTL/cortexm0ds_logic.v(19161)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5314|_al_u5313  (
    .a({_al_u5312_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({_al_u5313_o,_al_u5067_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5opw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 ,_al_u5313_o}));
  // ../RTL/cortexm0ds_logic.v(18172)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5315|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n48061}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,open_n48062}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5315_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 }),
    .q({open_n48083,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 }));  // ../RTL/cortexm0ds_logic.v(18172)
  // ../RTL/cortexm0ds_logic.v(18190)
  EG_PHY_LSLICE #(
    //.LUTF0("(D@(B*~(~C*A)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(D@(B*~(~C*A)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011101111000100),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0011101111000100),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5316|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 ,_al_u4219_o}),
    .b({_al_u5315_o,_al_u5620_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,_al_u5523_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 }),
    .mi({open_n48087,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 }),
    .f({_al_u5316_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[5]_i1[5]_o_lutinv }),
    .q({open_n48103,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Npaax6 }));  // ../RTL/cortexm0ds_logic.v(18190)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5319|_al_u5318  (
    .a({_al_u5311_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({_al_u5316_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5317_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc5bx6 }),
    .d({_al_u5318_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 }),
    .f({_al_u5319_o,_al_u5318_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u531|_al_u1676  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ,_al_u1676_o}));
  // ../RTL/cortexm0ds_logic.v(19887)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5321|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6_reg  (
    .b({_al_u5020_o,_al_u5053_o}),
    .c({_al_u5320_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }),
    .clk(XTAL1_wire),
    .d({_al_u5310_o,_al_u5321_o}),
    .f({_al_u5321_o,open_n48168}),
    .q({open_n48172,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ceabx6 }));  // ../RTL/cortexm0ds_logic.v(19887)
  // ../RTL/cortexm0ds_logic.v(20150)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5323|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5323_o,open_n48186}),
    .q({open_n48190,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 }));  // ../RTL/cortexm0ds_logic.v(20150)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*A*~(D*C))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"))
    \_al_u5324|_al_u6757  (
    .a({_al_u5323_o,open_n48191}),
    .b({_al_u5260_o,_al_u5260_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rzciu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtjow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }),
    .f({_al_u5324_o,_al_u6757_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5326|_al_u5325  (
    .a({_al_u5324_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({_al_u5325_o,_al_u5067_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oyhbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 ,_al_u5325_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5327|_al_u613  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .c({_al_u5275_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .d({_al_u374_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .f({_al_u5327_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 }));
  // ../RTL/cortexm0ds_logic.v(18595)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(D*~(C*B)))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("~(~A*~(D*~(C*B)))"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111110101010),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1011111110101010),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5328|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6_reg  (
    .a({open_n48258,_al_u1779_o}),
    .b({_al_u5327_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5328_o,open_n48276}),
    .q({open_n48280,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thiax6 }));  // ../RTL/cortexm0ds_logic.v(18595)
  // ../RTL/cortexm0ds_logic.v(18006)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5329|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6_reg  (
    .a({open_n48281,_al_u926_o}),
    .b({open_n48282,_al_u927_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .mi({open_n48293,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .f({_al_u5329_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 }),
    .q({open_n48298,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bt2qw6 }));  // ../RTL/cortexm0ds_logic.v(18006)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5332|_al_u5331  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 ,open_n48299}),
    .b({_al_u5328_o,_al_u1385_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] }),
    .d({_al_u5331_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .f({_al_u5332_o,_al_u5331_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5337|_al_u5334  (
    .a({_al_u5333_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({_al_u5334_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5335_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5yax6 }),
    .d({_al_u5336_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 }),
    .f({_al_u5337_o,_al_u5334_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D)*~(B)*~(C)+D*B*~(C)+~(D)*~(B)*C+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*C*~B*A)"),
    .INIT_LUT0(16'b1100110011110011),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"))
    \_al_u5339|_al_u5338  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ,open_n48344}),
    .b({_al_u5338_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .f({_al_u5339_o,_al_u5338_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u533|_al_u509  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .f({_al_u533_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~B*~(~D*C*A))"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~B*~(~D*C*A))"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0011001100010011),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0011001100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5340|_al_u5291  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 }),
    .b({_al_u5339_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .f({_al_u5340_o,_al_u5291_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5341|_al_u5647  (
    .b({open_n48415,_al_u5275_o}),
    .c({_al_u5275_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 }),
    .f({_al_u5341_o,_al_u5647_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~B*A*~(D*C))"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"))
    \_al_u5343|_al_u5342  (
    .a({_al_u5340_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv }),
    .b({_al_u5341_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ilwiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+~(A)*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    //.LUT1("(~C*B*~(~D*~A))"),
    .INIT_LUT0(16'b1110011000000000),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"))
    \_al_u5345|_al_u5344  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H2qiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D43qw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .c({_al_u5344_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe7ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .f({_al_u5345_o,_al_u5344_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5346|_al_u506  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .d({_al_u5345_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .f({_al_u5346_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~D*C*B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000000010000000),
    .MODE("LOGIC"))
    \_al_u5347|_al_u5699  (
    .a({_al_u5332_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .b({_al_u5337_o,_al_u5693_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv ,_al_u5698_o}),
    .d({_al_u5346_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvpiu6_lutinv }),
    .f({_al_u5347_o,_al_u5699_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(D*~C)))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(A*~(B*~(D*~C)))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0010101000100010),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0010101000100010),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5349|_al_u5348  (
    .a({open_n48524,_al_u5020_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5347_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 ,_al_u4637_o}),
    .d({_al_u5348_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5349_o,_al_u5348_o}));
  // ../RTL/cortexm0ds_logic.v(18289)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5351|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,open_n48549}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ,open_n48550}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 }),
    .mi({open_n48554,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({_al_u5351_o,_al_u5644_o}),
    .q({open_n48570,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 }));  // ../RTL/cortexm0ds_logic.v(18289)
  // ../RTL/cortexm0ds_logic.v(18311)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(~C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101000111110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5353|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u4423_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 ,_al_u5791_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 ,_al_u5800_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 }),
    .mi({open_n48581,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({_al_u5353_o,_al_u5801_o}),
    .q({open_n48586,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tceax6 }));  // ../RTL/cortexm0ds_logic.v(18311)
  // ../RTL/cortexm0ds_logic.v(18175)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~(D@A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*B*~(D@A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000001000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1000000001000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5354|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kikhu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,_al_u5501_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 ,_al_u5510_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 }),
    .mi({open_n48590,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({_al_u5354_o,_al_u5511_o}),
    .q({open_n48606,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lx9ax6 }));  // ../RTL/cortexm0ds_logic.v(18175)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5355|_al_u5352  (
    .a({_al_u5352_o,open_n48607}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wzpiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .c({_al_u5353_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 }),
    .d({_al_u5354_o,_al_u5351_o}),
    .f({_al_u5355_o,_al_u5352_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5356|_al_u1385  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 }),
    .d({_al_u927_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv ,_al_u1385_o}));
  // ../RTL/cortexm0ds_logic.v(18205)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5357|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv ,open_n48656}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fm7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbfax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .mi({open_n48667,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5357_o,_al_u5395_o}),
    .q({open_n48671,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0bax6 }));  // ../RTL/cortexm0ds_logic.v(18205)
  // ../RTL/cortexm0ds_logic.v(18231)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111011101000101),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111011101000101),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5358|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ,_al_u5643_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,_al_u5644_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5358_o,open_n48689}),
    .q({open_n48693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkbax6 }));  // ../RTL/cortexm0ds_logic.v(18231)
  // ../RTL/cortexm0ds_logic.v(18151)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5359|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6_reg  (
    .b({_al_u5345_o,open_n48696}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5359_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .q({open_n48712,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vz8ax6 }));  // ../RTL/cortexm0ds_logic.v(18151)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u5360|_al_u5696  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nu5bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xrxax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 }),
    .f({_al_u5360_o,_al_u5696_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5361|_al_u5362  (
    .a({open_n48733,_al_u5357_o}),
    .b({_al_u5359_o,_al_u5361_o}),
    .c({_al_u5360_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .d({_al_u5358_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] }),
    .f({_al_u5361_o,_al_u5362_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u5363|_al_u5290  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .c({_al_u5338_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .d({_al_u5346_o,_al_u5275_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffqiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5364|_al_u5661  (
    .a({open_n48776,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({open_n48777,_al_u405_o}),
    .c({_al_u5260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6rpw6 }),
    .d({_al_u405_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 }),
    .f({_al_u5364_o,_al_u5661_o}));
  // ../RTL/cortexm0ds_logic.v(19908)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110001000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1101111110001000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5365|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5365_o,open_n48819}),
    .q({open_n48823,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 }));  // ../RTL/cortexm0ds_logic.v(19908)
  // ../RTL/cortexm0ds_logic.v(19065)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5368|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6_reg  (
    .a({_al_u5364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({_al_u5365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 }),
    .c({_al_u5366_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dooow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 }),
    .mi({open_n48834,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 ,_al_u5366_o}),
    .q({open_n48838,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I2zax6 }));  // ../RTL/cortexm0ds_logic.v(19065)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*~(D*~B)))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0010101000001010),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5369|_al_u5370  (
    .a({_al_u5355_o,_al_u5020_o}),
    .b({_al_u5362_o,_al_u4611_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ,_al_u5369_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5369_o,_al_u5370_o}));
  // ../RTL/cortexm0ds_logic.v(18098)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5371|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 }),
    .clk(XTAL1_wire),
    .d({_al_u5370_o,_al_u5371_o}),
    .f({_al_u5371_o,open_n48875}),
    .q({open_n48879,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg7ax6 }));  // ../RTL/cortexm0ds_logic.v(18098)
  // ../RTL/cortexm0ds_logic.v(18401)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5373|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,_al_u5812_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,_al_u5813_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 ,_al_u5759_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 }),
    .mi({open_n48883,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mq1iu6 ,_al_u5814_o}),
    .q({open_n48899,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K6gax6 }));  // ../RTL/cortexm0ds_logic.v(18401)
  // ../RTL/cortexm0ds_logic.v(18402)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5374|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,_al_u5730_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,_al_u5809_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 }),
    .mi({open_n48903,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu1iu6 ,_al_u5813_o}),
    .q({open_n48919,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H8gax6 }));  // ../RTL/cortexm0ds_logic.v(18402)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*~(D*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0100000011000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5376|_al_u5375  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uu1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5375_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usnpw6 }),
    .f({_al_u5376_o,_al_u5375_o}));
  // ../RTL/cortexm0ds_logic.v(18403)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5377|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mq1iu6 ,_al_u2150_o}),
    .b({_al_u5376_o,_al_u2272_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n48954,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .f({_al_u5377_o,_al_u2274_o}),
    .q({open_n48959,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 }));  // ../RTL/cortexm0ds_logic.v(18403)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C*B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(A*~(D*C*B))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b0010101010101010),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0010101010101010),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5378|_al_u5389  (
    .a({open_n48960,_al_u5020_o}),
    .b({_al_u1865_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,_al_u5378_o}),
    .d({_al_u5377_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 }),
    .f({_al_u5378_o,_al_u5389_o}));
  // ../RTL/cortexm0ds_logic.v(20219)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5379|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [31]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5379_o,open_n48998}),
    .q({open_n49002,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 }));  // ../RTL/cortexm0ds_logic.v(20219)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(C*~B*D)"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"))
    \_al_u537|_al_u534  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqwpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zm8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cvciu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5383|_al_u5381  (
    .a({open_n49025,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 }),
    .b({_al_u5381_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 }),
    .c({_al_u5382_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 }),
    .d({_al_u5380_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 }),
    .f({_al_u5383_o,_al_u5381_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5385|_al_u5384  (
    .a({open_n49046,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 }),
    .d({_al_u5384_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 }),
    .f({_al_u5385_o,_al_u5384_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5388|_al_u5387  (
    .a({_al_u5383_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .b({_al_u5385_o,_al_u3779_o}),
    .c({_al_u5386_o,_al_u5260_o}),
    .d({_al_u5387_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 ,_al_u5387_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u538|_al_u514  (
    .b({open_n49097,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0xiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hw8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xiu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }));
  // ../RTL/cortexm0ds_logic.v(17478)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5390|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6_reg  (
    .a({_al_u5389_o,open_n49122}),
    .b({_al_u5050_o,_al_u5053_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 ,_al_u5390_o}),
    .f({_al_u5390_o,open_n49137}),
    .q({open_n49141,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 }));  // ../RTL/cortexm0ds_logic.v(17478)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5392|_al_u5706  (
    .a({open_n49142,_al_u5392_o}),
    .b({open_n49143,_al_u5705_o}),
    .c({_al_u4368_o,_al_u3887_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E18iu6 ,_al_u3889_o}),
    .f({_al_u5392_o,_al_u5706_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5393|_al_u3162  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u5392_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1465 }));
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111001100),
    .INIT_LUT1(16'b1010001010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5394|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/wr_reg_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ,open_n49188}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq4iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5394_o,\u_cmsdk_mcu/HWRITE }),
    .q({open_n49204,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5397|_al_u5489  (
    .b({open_n49207,_al_u5399_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] }),
    .d({_al_u5396_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7],_al_u5489_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5398|_al_u5396  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 }),
    .d({_al_u5395_o,_al_u5395_o}),
    .f({_al_u5398_o,_al_u5396_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*A*~(~C*B))"),
    //.LUTF1("(C*B*~(~D*~A))"),
    //.LUTG0("(~D*A*~(~C*B))"),
    //.LUTG1("(C*B*~(~D*~A))"),
    .INIT_LUTF0(16'b0000000010100010),
    .INIT_LUTF1(16'b1100000010000000),
    .INIT_LUTG0(16'b0000000010100010),
    .INIT_LUTG1(16'b1100000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5401|_al_u5400  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ,_al_u5398_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7],_al_u5399_o}),
    .c({_al_u5400_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .d({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chkhu6 ,_al_u5400_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5403|_al_u5335  (
    .a({open_n49280,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({open_n49281,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 }),
    .d({_al_u5395_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 }),
    .f({_al_u5403_o,_al_u5335_o}));
  // ../RTL/cortexm0ds_logic.v(18220)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~C*~B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5404|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ,_al_u5403_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5403_o,_al_u5396_o}),
    .mi({open_n49307,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [3],_al_u5474_o}),
    .q({open_n49323,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 }));  // ../RTL/cortexm0ds_logic.v(18220)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(~D*~B)))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~A*~(C*~(~D*~B)))"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000010100010101),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000010100010101),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5405|_al_u5479  (
    .a({open_n49324,_al_u5396_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ,_al_u5398_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ,_al_u5403_o}),
    .d({_al_u5395_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ,_al_u5479_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b1100010000000100),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1100010000000100),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5406|_al_u5503  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ,_al_u4225_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ,_al_u5399_o}),
    .d({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufkhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjkhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5407|_al_u7156  (
    .a({open_n49373,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] }),
    .d({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [3]}),
    .f({_al_u5407_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkfow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(D*B*~(~C*~A))"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(D*B*~(~C*~A))"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b1100100000000000),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b1100100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5408|_al_u5409  (
    .a({_al_u5398_o,open_n49398}),
    .b({_al_u5403_o,_al_u5408_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ,_al_u5399_o}),
    .d({_al_u5407_o,_al_u4231_o}),
    .f({_al_u5408_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5410|_al_u5430  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7bax6 ,_al_u5403_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 }),
    .d({_al_u5395_o,_al_u5398_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ,_al_u5430_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~B*D))"),
    //.LUT1("(C*B*~D)"),
    .INIT_LUT0(16'b0000110000001111),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"))
    \_al_u5413|_al_u5412  (
    .b({_al_u5403_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] }),
    .c({_al_u5412_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 }),
    .d({_al_u5411_o,_al_u5399_o}),
    .f({_al_u5413_o,_al_u5412_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u5414|_al_u5535  (
    .b({_al_u5413_o,_al_u5534_o}),
    .c({_al_u5399_o,_al_u5523_o}),
    .d({_al_u4141_o,_al_u4141_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(~D*A))"),
    //.LUTF1("(~(~C*B)*~(D*~A))"),
    //.LUTG0("(~(~C*B)*~(~D*A))"),
    //.LUTG1("(~(~C*B)*~(D*~A))"),
    .INIT_LUTF0(16'b1111001101010001),
    .INIT_LUTF1(16'b1010001011110011),
    .INIT_LUTG0(16'b1111001101010001),
    .INIT_LUTG1(16'b1010001011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5415|_al_u5473  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alkhu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 }),
    .f({_al_u5415_o,_al_u5473_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*C))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u5418|_al_u5417  (
    .a({open_n49517,_al_u5416_o}),
    .b({_al_u5417_o,_al_u5396_o}),
    .c({_al_u5399_o,_al_u5399_o}),
    .d({_al_u4106_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqkhu6 ,_al_u5417_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(D*~(C@B))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5419|_al_u5478  (
    .a({open_n49538,_al_u5470_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqkhu6 ,_al_u5473_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fo9ax6 ,_al_u5476_o}),
    .d({_al_u5415_o,_al_u5477_o}),
    .f({_al_u5419_o,_al_u5478_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5420|_al_u5399  (
    .c({_al_u5403_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 }),
    .d({_al_u5396_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 }),
    .f({_al_u5420_o,_al_u5399_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5421|_al_u5422  (
    .a({open_n49591,_al_u3889_o}),
    .b({open_n49592,_al_u5421_o}),
    .c({_al_u5411_o,_al_u5399_o}),
    .d({_al_u5420_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] }),
    .f({_al_u5421_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5424|_al_u5283  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 }),
    .f({_al_u5424_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tsriu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u5426|_al_u5425  (
    .b({_al_u5425_o,_al_u5399_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] }),
    .d({_al_u5411_o,_al_u5396_o}),
    .f({_al_u5426_o,_al_u5425_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .INIT_LUT0(16'b1100010000000100),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"))
    \_al_u5428|_al_u5423  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 ,_al_u4121_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nvkbx6 [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bq9ax6 ,_al_u5399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] }),
    .f({_al_u5428_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yokhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5429|_al_u5446  (
    .b({_al_u5424_o,open_n49685}),
    .c({_al_u5428_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J59ax6 }),
    .d({_al_u5419_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uilhu6 }),
    .f({_al_u5429_o,_al_u5446_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5431|_al_u5432  (
    .a({open_n49710,_al_u4191_o}),
    .b({open_n49711,_al_u5431_o}),
    .c({_al_u5396_o,_al_u5399_o}),
    .d({_al_u5430_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] }),
    .f({_al_u5431_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5433|_al_u5411  (
    .b({_al_u5395_o,_al_u5395_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv }),
    .f({_al_u5433_o,_al_u5411_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5434|_al_u5460  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ,_al_u5396_o}),
    .d({_al_u5403_o,_al_u5416_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv ,_al_u5460_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5435|_al_u5436  (
    .a({open_n49782,_al_u4081_o}),
    .b({open_n49783,_al_u5435_o}),
    .c({_al_u5396_o,_al_u5399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] }),
    .f({_al_u5435_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7lhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5439|_al_u5438  (
    .b({_al_u5403_o,_al_u5399_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] }),
    .d({_al_u5438_o,_al_u5396_o}),
    .f({_al_u5439_o,_al_u5438_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u543|_al_u284  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ,open_n49830}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ,open_n49831}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .f({_al_u543_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [1]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"))
    \_al_u5441|_al_u5440  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 ,open_n49852}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lclhu6 ,_al_u5439_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G79ax6 ,_al_u5399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 ,_al_u4126_o}),
    .f({_al_u5441_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 }));
  // ../RTL/cortexm0ds_logic.v(18221)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~D*~C*B))"),
    //.LUTF1("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG0("(~A*~(~D*~C*B))"),
    //.LUTG1("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010101010001),
    .INIT_LUTF1(16'b0011000100000001),
    .INIT_LUTG0(16'b0101010101010001),
    .INIT_LUTG1(16'b0011000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5443|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6_reg  (
    .a({_al_u4061_o,_al_u5396_o}),
    .b({_al_u5442_o,_al_u5398_o}),
    .c({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 }),
    .mi({open_n49876,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2lhu6 ,_al_u5442_o}),
    .q({open_n49892,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9bax6 }));  // ../RTL/cortexm0ds_logic.v(18221)
  // ../RTL/cortexm0ds_logic.v(19933)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("~(C@D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("~(C@D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111000000001111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5444|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6_reg  (
    .a({open_n49893,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({open_n49894,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2lhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 }),
    .mi({open_n49898,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .f({_al_u5444_o,_al_u6665_o}),
    .q({open_n49914,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjbbx6 }));  // ../RTL/cortexm0ds_logic.v(19933)
  // ../RTL/cortexm0ds_logic.v(19987)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C@B))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100001100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5445|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6_reg  (
    .a({_al_u5429_o,open_n49915}),
    .b({_al_u5437_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G7lhu6 }),
    .c({_al_u5441_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5444_o,_al_u5433_o}),
    .mi({open_n49926,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .f({_al_u5445_o,_al_u5437_o}),
    .q({open_n49931,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M4ebx6 }));  // ../RTL/cortexm0ds_logic.v(19987)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~D*~C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(~D*~C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0011001100110001),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011001100110001),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5447|_al_u5416  (
    .a({open_n49932,_al_u5398_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ,_al_u5403_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 }),
    .d({_al_u5398_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5bax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ,_al_u5416_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5448|_al_u5467  (
    .c({_al_u5403_o,_al_u5396_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv }),
    .f({_al_u5448_o,_al_u5467_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5449|_al_u5450  (
    .a({open_n49981,_al_u4096_o}),
    .b({open_n49982,_al_u5449_o}),
    .c({_al_u5396_o,_al_u5399_o}),
    .d({_al_u5448_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] }),
    .f({_al_u5449_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u544|_al_u280  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ,open_n50003}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ,open_n50004}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .f({_al_u544_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D@A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(C*~B)*~(D@A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1000101001000101),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1000101001000101),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5451|_al_u5457  (
    .a({open_n50025,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eukhu6 }),
    .b({open_n50026,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sdlhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv8bx6 }),
    .f({_al_u5451_o,_al_u5457_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUT1("~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    .INIT_LUT0(16'b0011111100001100),
    .INIT_LUT1(16'b0011111100001100),
    .MODE("LOGIC"))
    \_al_u5452|_al_u5598  (
    .b({_al_u5399_o,_al_u5523_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] }),
    .d({_al_u3887_o,_al_u3887_o}),
    .f({_al_u5452_o,_al_u5598_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5455|_al_u5454  (
    .b({_al_u5398_o,_al_u5399_o}),
    .c({_al_u5403_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] }),
    .d({_al_u5454_o,_al_u5396_o}),
    .f({_al_u5455_o,_al_u5454_o}));
  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5456|u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/reg0_b9  (
    .b({_al_u5455_o,_al_u4116_o}),
    .c({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/trans_valid ),
    .clk(XTAL1_wire),
    .d({_al_u4116_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eukhu6 ,\u_cmsdk_mcu/HADDR [11]}),
    .q({open_n50121,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_system_rom_table/haddr_reg [9]}));  // ../RTL/cmsdk_ahb_cs_rom_table.v(161)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u5458|_al_u5459  (
    .a({open_n50122,_al_u4101_o}),
    .b({_al_u5398_o,_al_u5458_o}),
    .c({_al_u5403_o,_al_u5399_o}),
    .d({_al_u5396_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] }),
    .f({_al_u5458_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 }));
  // ../RTL/cortexm0ds_logic.v(18571)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(C*~(B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1100111100001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u545|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6_reg  (
    .b({_al_u544_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 }),
    .clk(XTAL1_wire),
    .d({_al_u543_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n3685 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 ,open_n50158}),
    .q({open_n50162,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daiax6 }));  // ../RTL/cortexm0ds_logic.v(18571)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0011000100000001),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0011000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5461|_al_u7210  (
    .a({_al_u4184_o,_al_u4289_o}),
    .b({_al_u5460_o,_al_u4290_o}),
    .c({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [23]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqcow6 }));
  // ../RTL/cortexm0ds_logic.v(19962)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(~(~C*B)*~(D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b1010001011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5462|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zelhu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 }),
    .mi({open_n50197,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .f({_al_u5462_o,_al_u5484_o}),
    .q({open_n50202,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Itcbx6 }));  // ../RTL/cortexm0ds_logic.v(19962)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5463|_al_u5464  (
    .a({open_n50203,_al_u4086_o}),
    .b({_al_u5396_o,_al_u5463_o}),
    .c({_al_u5403_o,_al_u5399_o}),
    .d({_al_u5411_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] }),
    .f({_al_u5463_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"))
    \_al_u5465|_al_u5470  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eblhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O8lhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D99ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 }),
    .f({_al_u5465_o,_al_u5470_o}));
  // ../RTL/cortexm0ds_logic.v(18399)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*(D@C))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~B*~A*(D@C))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100010000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000100010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5466|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6_reg  (
    .a({_al_u5453_o,_al_u5446_o}),
    .b({_al_u5457_o,_al_u5451_o}),
    .c({_al_u5462_o,_al_u5452_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5465_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 }),
    .mi({open_n50251,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .f({_al_u5466_o,_al_u5453_o}),
    .q({open_n50267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2gax6 }));  // ../RTL/cortexm0ds_logic.v(18399)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~(~D*A))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(C*~B*~(~D*A))"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0011000000010000),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5468|_al_u5469  (
    .a({open_n50268,_al_u4066_o}),
    .b({_al_u5399_o,_al_u5467_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ,_al_u5468_o}),
    .d({_al_u5420_o,_al_u5399_o}),
    .f({_al_u5468_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*C))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u5472|_al_u5471  (
    .a({open_n50293,_al_u5448_o}),
    .b({_al_u5471_o,_al_u5396_o}),
    .c({_al_u5399_o,_al_u5399_o}),
    .d({_al_u4111_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 ,_al_u5471_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"))
    \_al_u5476|_al_u5427  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 ,open_n50314}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 ,_al_u5426_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ,_al_u5399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 ,_al_u4131_o}),
    .f({_al_u5476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cykhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0011000100000001),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0011000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5480|_al_u7080  (
    .a({_al_u4076_o,_al_u4289_o}),
    .b({_al_u5479_o,_al_u4290_o}),
    .c({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [19]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 ,_al_u7080_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(~D*C))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(B*~A*~(~D*C))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0100010000000100),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5483|_al_u5482  (
    .a({open_n50359,_al_u5430_o}),
    .b({_al_u5482_o,_al_u5396_o}),
    .c({_al_u5399_o,_al_u5399_o}),
    .d({_al_u4237_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 ,_al_u5482_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5487|_al_u5486  (
    .a({_al_u5481_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 }),
    .b({_al_u5484_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwkhu6 }),
    .c({_al_u5485_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 }),
    .d({_al_u5486_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 }),
    .f({_al_u5487_o,_al_u5486_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~(D@A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*B*~(D@A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1000000001000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000000001000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5488|_al_u5513  (
    .a({_al_u5445_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufkhu6 }),
    .b({_al_u5466_o,_al_u5488_o}),
    .c({_al_u5478_o,_al_u5511_o}),
    .d({_al_u5487_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttmhu6 }),
    .f({_al_u5488_o,_al_u5513_o}));
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*B*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1100000001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5490|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b5  (
    .a({_al_u4423_o,open_n50432}),
    .b({_al_u5489_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6018_lutinv ,_al_u4423_o}),
    .clk(XTAL1_wire),
    .d({_al_u5399_o,\u_cmsdk_mcu/HADDR [5]}),
    .mi({open_n50444,\u_cmsdk_mcu/HADDR [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kikhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bg9iu6 }),
    .q({open_n50448,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cortexm0ds_logic.v(18166)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C@D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5492|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6_reg  (
    .a({open_n50449,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({open_n50450,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzkhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 }),
    .mi({open_n50454,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[15]_i1[15]_o_lutinv ,_al_u6699_o}),
    .q({open_n50470,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rg9ax6 }));  // ../RTL/cortexm0ds_logic.v(18166)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~C*~B*~D)"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5493|_al_u5494  (
    .a({open_n50471,_al_u3885_o}),
    .b({_al_u5403_o,_al_u5493_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6021_lutinv ,_al_u5399_o}),
    .d({_al_u5396_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] }),
    .f({_al_u5493_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhlhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5495|_al_u5496  (
    .a({open_n50496,_al_u4197_o}),
    .b({_al_u5398_o,_al_u5495_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ,_al_u5399_o}),
    .d({_al_u5420_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] }),
    .f({_al_u5495_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gglhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u5498|_al_u5475  (
    .a({open_n50521,_al_u4071_o}),
    .b({_al_u5399_o,_al_u5474_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ,_al_u5399_o}),
    .d({_al_u5474_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] }),
    .f({_al_u5498_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u5499|_al_u5500  (
    .b({_al_u5396_o,_al_u5499_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ,_al_u5399_o}),
    .d({_al_u5498_o,_al_u4056_o}),
    .f({_al_u5499_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0lhu6 }));
  // ../RTL/cortexm0ds_logic.v(18165)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*~A*~(D@C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0100000000000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5501|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[15]_i1[15]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u5497_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0lhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 }),
    .mi({open_n50574,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .f({_al_u5501_o,_al_u6677_o}),
    .q({open_n50579,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ue9ax6 }));  // ../RTL/cortexm0ds_logic.v(18165)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0011000100000001),
    .MODE("LOGIC"))
    \_al_u5502|_al_u7087  (
    .a({_al_u4091_o,_al_u4289_o}),
    .b({_al_u5420_o,_al_u4290_o}),
    .c({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [22]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9lhu6 ,_al_u7087_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(~D*C))"),
    //.LUTF1("(D@(B*~(~C*A)))"),
    //.LUTG0("(B*A*~(~D*C))"),
    //.LUTG1("(D@(B*~(~C*A)))"),
    .INIT_LUTF0(16'b1000100000001000),
    .INIT_LUTF1(16'b0011101111000100),
    .INIT_LUTG0(16'b1000100000001000),
    .INIT_LUTG1(16'b0011101111000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5506|_al_u5505  (
    .a({_al_u4219_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6006_lutinv }),
    .b({_al_u5505_o,_al_u5396_o}),
    .c({_al_u5399_o,_al_u5399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xr9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[5]_i1[5]_o_lutinv ,_al_u5505_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*C))"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u5507|_al_u5508  (
    .a({open_n50624,_al_u5507_o}),
    .b({_al_u5403_o,_al_u5396_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n6023_lutinv ,_al_u5399_o}),
    .d({_al_u5398_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] }),
    .f({_al_u5507_o,_al_u5508_o}));
  // ../RTL/cortexm0ds_logic.v(18168)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D@(B*~(~C*A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011101111000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5509|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6_reg  (
    .a({_al_u4035_o,open_n50645}),
    .b({_al_u5508_o,open_n50646}),
    .c({_al_u5399_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .mi({open_n50657,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[12]_i1[12]_o_lutinv ,_al_u2085_o}),
    .q({open_n50662,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 }));  // ../RTL/cortexm0ds_logic.v(18168)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5510|_al_u2039  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[5]_i1[5]_o_lutinv ,open_n50665}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[12]_i1[12]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G30iu6 }),
    .d({_al_u5504_o,_al_u2038_o}),
    .f({_al_u5510_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 }));
  // ../RTL/cortexm0ds_logic.v(18159)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5512|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6_reg  (
    .a({open_n50690,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 }),
    .b({open_n50691,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 }),
    .mi({open_n50702,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttmhu6 ,_al_u5655_o}),
    .q({open_n50707,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N39ax6 }));  // ../RTL/cortexm0ds_logic.v(18159)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(C*~B*~(~D*~A))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0011000000100000),
    .MODE("LOGIC"))
    \_al_u5515|_al_u5514  (
    .a({_al_u5394_o,_al_u5399_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[1]_i1[1]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 }),
    .c({_al_u5513_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 }),
    .d({_al_u5514_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u5515_o,_al_u5514_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5516|_al_u5638  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv }),
    .f({_al_u5516_o,_al_u5638_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1010001010000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1010001010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5518|_al_u5523  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xipiu6 ,open_n50752}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnpiu6 ,open_n50753}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 }),
    .f({_al_u5518_o,_al_u5523_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5522|_al_u5520  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 }),
    .d({_al_u5519_o,_al_u5519_o}),
    .f({_al_u5522_o,_al_u5520_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*A*~(~D*B))"),
    //.LUT1("(C*B*~(~D*~A))"),
    .INIT_LUT0(16'b0000101000000010),
    .INIT_LUT1(16'b1100000010000000),
    .MODE("LOGIC"))
    \_al_u5525|_al_u5524  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 ,_al_u5522_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7],_al_u5523_o}),
    .c({_al_u5524_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 }),
    .d({_al_u5523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhhu6 ,_al_u5524_o}));
  // ../RTL/cortexm0ds_logic.v(18194)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(A@(D*~(~C*~B)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0101011010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5526|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxhhu6 ,open_n50826}),
    .b({_al_u1888_o,open_n50827}),
    .c({_al_u5523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8ipw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[1]_i1[1]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .q({open_n50844,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 }));  // ../RTL/cortexm0ds_logic.v(18194)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5527|_al_u5559  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 ,_al_u5522_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 }),
    .d({_al_u5522_o,_al_u5520_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [3],_al_u5559_o}));
  // ../RTL/cortexm0ds_logic.v(20254)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*A*~(D*C))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~B*A*~(D*C))"),
    //.LUTG1("(~C*~B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000100010),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5528|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6_reg  (
    .a({open_n50871,_al_u5519_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5519_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 }),
    .mi({open_n50875,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv }),
    .q({open_n50891,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 }));  // ../RTL/cortexm0ds_logic.v(20254)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b1100010000000100),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1100010000000100),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5529|_al_u5611  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/My0iu6 ,_al_u4225_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ,_al_u5523_o}),
    .d({_al_u5523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwhhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0ihu6 }));
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u552|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b9  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [8],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [13]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u552_o,open_n50934}),
    .q({open_n50938,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [9]}));  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u5531|_al_u5605  (
    .b({_al_u5519_o,_al_u5532_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ,_al_u5520_o}),
    .f({_al_u5531_o,_al_u5605_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5532|_al_u5521  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 }),
    .d({_al_u5519_o,_al_u5520_o}),
    .f({_al_u5532_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~B*D))"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~C*~(~B*D))"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0000110000001111),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000110000001111),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5534|_al_u5533  (
    .b({_al_u5532_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] }),
    .c({_al_u5533_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 }),
    .d({_al_u5531_o,_al_u5523_o}),
    .f({_al_u5534_o,_al_u5533_o}));
  // ../RTL/cortexm0ds_logic.v(18226)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(C*A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b1000000010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5537|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6_reg  (
    .a({_al_u5532_o,open_n51011}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 }),
    .c({_al_u5536_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ,_al_u5523_o}),
    .mi({open_n51022,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .f({_al_u5537_o,_al_u5536_o}),
    .q({open_n51027,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 }));  // ../RTL/cortexm0ds_logic.v(18226)
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u553|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [3],open_n51028}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [10]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u553_o,open_n51045}),
    .q({open_n51049,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [6]}));  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~A*~(~D*B))"),
    //.LUTF1("(A*~(~C*~(~D*B)))"),
    //.LUTG0("(~C*~A*~(~D*B))"),
    //.LUTG1("(A*~(~C*~(~D*B)))"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b1010000010101000),
    .INIT_LUTG0(16'b0000010100000001),
    .INIT_LUTG1(16'b1010000010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5540|_al_u5588  (
    .a({_al_u5520_o,_al_u5520_o}),
    .b({_al_u5522_o,_al_u5522_o}),
    .c({_al_u5532_o,_al_u5532_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [9],_al_u5588_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5541|_al_u5594  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ,open_n51076}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv }),
    .d({_al_u5519_o,_al_u5520_o}),
    .f({_al_u5541_o,_al_u5594_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(C*B*~(~D*A))"),
    //.LUTG0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(C*B*~(~D*A))"),
    .INIT_LUTF0(16'b1100010000000100),
    .INIT_LUTF1(16'b1100000001000000),
    .INIT_LUTG0(16'b1100010000000100),
    .INIT_LUTG1(16'b1100000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5543|_al_u5566  (
    .a({_al_u4106_o,_al_u4237_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [9]}),
    .c({_al_u5542_o,_al_u5523_o}),
    .d({_al_u5523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S6ihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5546|_al_u5198  (
    .b({open_n51127,_al_u1385_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] }),
    .d({_al_u5523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .f({_al_u5546_o,_al_u5198_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(~D*~(~A*~(C*B)))"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(~D*~(~A*~(C*B)))"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b0000000011101010),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b0000000011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5547|_al_u5548  (
    .a({_al_u5520_o,open_n51148}),
    .b({_al_u5532_o,_al_u5547_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ,_al_u5523_o}),
    .d({_al_u5546_o,_al_u4066_o}),
    .f({_al_u5547_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(~(C*~B)*~(~D*A))"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(~(C*~B)*~(~D*A))"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b1100111101000101),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b1100111101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5549|_al_u5538  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 ,open_n51173}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 ,_al_u5537_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ,_al_u4231_o}),
    .f({_al_u5549_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 }));
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u554|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [13],open_n51198}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u554_o,open_n51215}),
    .q({open_n51219,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [2]}));  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~A*~(~D*~C*B))"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~A*~(~D*~C*B))"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b0101010101010001),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5550|_al_u5551  (
    .a({_al_u5520_o,_al_u4061_o}),
    .b({_al_u5522_o,_al_u5550_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] }),
    .f({_al_u5550_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miihu6 }));
  // ../RTL/cortexm0ds_logic.v(19934)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5552|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6_reg  (
    .a({_al_u5544_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .b({_al_u5549_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pbbbx6 }),
    .mi({open_n51254,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .f({_al_u5552_o,_al_u6663_o}),
    .q({open_n51259,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlbbx6 }));  // ../RTL/cortexm0ds_logic.v(19934)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u5554|_al_u5553  (
    .b({_al_u5553_o,_al_u5523_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] }),
    .d({_al_u5531_o,_al_u5520_o}),
    .f({_al_u5554_o,_al_u5553_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5556|_al_u5555  (
    .b({open_n51284,_al_u5554_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 ,_al_u4131_o}),
    .f({_al_u5556_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u555|_al_u618  (
    .b({_al_u553_o,open_n51311}),
    .c({_al_u554_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated }),
    .d({_al_u552_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i }),
    .f({_al_u555_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~A*~(B*~(D*~C)))"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0001010100010001),
    .MODE("LOGIC"))
    \_al_u5562|_al_u5563  (
    .a({_al_u5520_o,_al_u4076_o}),
    .b({_al_u5532_o,_al_u5562_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] }),
    .f({_al_u5562_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5565|_al_u5582  (
    .a({_al_u5552_o,_al_u5573_o}),
    .b({_al_u5558_o,_al_u5577_o}),
    .c({_al_u5561_o,_al_u5580_o}),
    .d({_al_u5564_o,_al_u5581_o}),
    .f({_al_u5565_o,_al_u5582_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5568|_al_u5567  (
    .b({_al_u5532_o,_al_u5523_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] }),
    .d({_al_u5567_o,_al_u5520_o}),
    .f({_al_u5568_o,_al_u5567_o}));
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u556|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [1],open_n51402}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [5]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u556_o,open_n51415}),
    .q({open_n51419,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [1]}));  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cortexm0ds_logic.v(18185)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(~C*B)*~(D*~A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(~C*B)*~(D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010001011110011),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010001011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5570|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 ,open_n51420}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 ,open_n51421}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .mi({open_n51425,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .f({_al_u5570_o,_al_u2107_o}),
    .q({open_n51441,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 }));  // ../RTL/cortexm0ds_logic.v(18185)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u5571|_al_u5572  (
    .a({open_n51442,_al_u4096_o}),
    .b({_al_u5532_o,_al_u5571_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ,_al_u5523_o}),
    .d({_al_u5520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] }),
    .f({_al_u5571_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guihu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C@B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"))
    \_al_u5573|_al_u5098  (
    .a({open_n51463,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Guihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cccbx6 }),
    .d({_al_u5570_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 }),
    .f({_al_u5573_o,_al_u5098_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5575|_al_u5574  (
    .b({_al_u5532_o,_al_u5523_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] }),
    .d({_al_u5574_o,_al_u5520_o}),
    .f({_al_u5575_o,_al_u5574_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(~B*~(C*~D))"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0011001100000011),
    .MODE("LOGIC"))
    \_al_u5578|_al_u5579  (
    .a({open_n51510,_al_u4086_o}),
    .b({_al_u5520_o,_al_u5578_o}),
    .c({_al_u5532_o,_al_u5523_o}),
    .d({_al_u5531_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] }),
    .f({_al_u5578_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 }));
  // ../RTL/cortexm0ds_logic.v(20014)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(~D*A))"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110001010100),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5580|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apihu6 ,_al_u5598_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 }),
    .mi({open_n51541,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .f({_al_u5580_o,_al_u5599_o}),
    .q({open_n51546,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlfbx6 }));  // ../RTL/cortexm0ds_logic.v(20014)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5583|_al_u5569  (
    .b({open_n51549,_al_u5568_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 ,_al_u4126_o}),
    .f({_al_u5583_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdihu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5585|_al_u5617  (
    .a({open_n51574,_al_u4091_o}),
    .b({open_n51575,_al_u5584_o}),
    .c({_al_u5584_o,_al_u5523_o}),
    .d({_al_u5531_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] }),
    .f({_al_u5585_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqihu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u5587|_al_u5586  (
    .a({open_n51596,_al_u3889_o}),
    .b({open_n51597,_al_u5585_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] }),
    .f({_al_u5587_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~B*~A*~(D@C))"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~B*~A*~(D@C))"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b0001000000000001),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b0001000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5590|_al_u5589  (
    .a({_al_u5583_o,_al_u4191_o}),
    .b({_al_u5587_o,_al_u5588_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysihu6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] }),
    .f({_al_u5590_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysihu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5591|_al_u5584  (
    .c({_al_u5532_o,_al_u5532_o}),
    .d({_al_u5522_o,_al_u5520_o}),
    .f({_al_u5591_o,_al_u5584_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5595|_al_u5596  (
    .a({open_n51670,_al_u4197_o}),
    .b({open_n51671,_al_u5595_o}),
    .c({_al_u5594_o,_al_u5523_o}),
    .d({_al_u5591_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] }),
    .f({_al_u5595_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwihu6 }));
  // ../RTL/cmsdk_apb_uart.v(476)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C@D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111100001010),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b1101111100001010),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u559|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_txd_reg  (
    .a({open_n51692,_al_u379_o}),
    .b({open_n51693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]}),
    .c({uart0_txd_pad,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_reg_txd ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_txd ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_reg_txd ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/nxt_txd }),
    .q({open_n51713,uart0_txd_pad}));  // ../RTL/cmsdk_apb_uart.v(476)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5600|_al_u5542  (
    .b({open_n51716,_al_u5523_o}),
    .c({_al_u5541_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] }),
    .d({_al_u5520_o,_al_u5541_o}),
    .f({_al_u5600_o,_al_u5542_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(~D*C))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0001000100000001),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u5602|_al_u5601  (
    .a({open_n51741,_al_u5588_o}),
    .b({_al_u5601_o,_al_u5600_o}),
    .c({_al_u5523_o,_al_u5523_o}),
    .d({_al_u4184_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qrihu6 ,_al_u5601_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(B*A*~(D@C))"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5607|_al_u5606  (
    .a({_al_u5603_o,_al_u3885_o}),
    .b({_al_u5604_o,_al_u5605_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyihu6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tchbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] }),
    .f({_al_u5607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyihu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(D@A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1000000001000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5608|_al_u5635  (
    .a({_al_u5565_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwhhu6 }),
    .b({_al_u5582_o,_al_u5608_o}),
    .c({_al_u5597_o,_al_u5633_o}),
    .d({_al_u5607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbkhu6 }),
    .f({_al_u5608_o,_al_u5635_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b1100010000000100),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1100010000000100),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5609|_al_u5557  (
    .a({open_n51806,_al_u4121_o}),
    .b({_al_u5523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntkbx6 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] }),
    .f({_al_u5609_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5ihu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5612|_al_u5336  (
    .a({open_n51831,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .b({open_n51832,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ftaax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E0ihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[3]_i1[3]_o_lutinv ,_al_u5336_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG0("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT_LUTF0(16'b1100010000000100),
    .INIT_LUTF1(16'b1100010000000100),
    .INIT_LUTG0(16'b1100010000000100),
    .INIT_LUTG1(16'b1100010000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5613|_al_u5491  (
    .a({_al_u4136_o,_al_u4136_o}),
    .b({_al_u5520_o,_al_u5396_o}),
    .c({_al_u5523_o,_al_u5399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzkhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~B*~A*~(~D*C))"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~B*~A*~(~D*C))"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b0001000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5614|_al_u5560  (
    .a({_al_u5594_o,_al_u4071_o}),
    .b({_al_u5559_o,_al_u5559_o}),
    .c({_al_u5523_o,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] }),
    .f({_al_u5614_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 }));
  // ../RTL/cortexm0ds_logic.v(18184)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~(C@D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~(C@D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011000000000011),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5616|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[16]_i1[16]_o_lutinv ,open_n51907}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .mi({open_n51911,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .f({_al_u5616_o,_al_u2151_o}),
    .q({open_n51927,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 }));  // ../RTL/cortexm0ds_logic.v(18184)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5620|_al_u5619  (
    .b({_al_u5532_o,_al_u5523_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] }),
    .d({_al_u5619_o,_al_u5520_o}),
    .f({_al_u5620_o,_al_u5619_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u5623|_al_u5622  (
    .b({_al_u5622_o,_al_u5523_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5997_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] }),
    .d({_al_u5591_o,_al_u5520_o}),
    .f({_al_u5623_o,_al_u5622_o}));
  // ../RTL/cortexm0ds_logic.v(18186)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(D@(B*~(~C*A)))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(D@(B*~(~C*A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0011101111000100),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0011101111000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5624|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6_reg  (
    .a({_al_u4035_o,open_n51972}),
    .b({_al_u5623_o,open_n51973}),
    .c({_al_u5523_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .mi({open_n51977,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[12]_i1[12]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 }),
    .q({open_n51993,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 }));  // ../RTL/cortexm0ds_logic.v(18186)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5625|_al_u5643  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[12]_i1[12]_o_lutinv ,_al_u5637_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[5]_i1[5]_o_lutinv ,_al_u5515_o}),
    .f({_al_u5625_o,_al_u5643_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(~D*C))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~A*~(~D*C))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0100010000000100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0100010000000100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5626|_al_u5592  (
    .a({open_n52018,_al_u5591_o}),
    .b({open_n52019,_al_u5520_o}),
    .c({_al_u5520_o,_al_u5523_o}),
    .d({_al_u5591_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] }),
    .f({_al_u5626_o,_al_u5592_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0011000100000001),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u5628|_al_u5627  (
    .a({open_n52044,_al_u4101_o}),
    .b({open_n52045,_al_u5626_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvcbx6 ,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[27]_i1[27]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovihu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~B*(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0011000100000001),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0011000100000001),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5629|_al_u5630  (
    .a({open_n52066,_al_u4081_o}),
    .b({_al_u5532_o,_al_u5629_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv ,_al_u5523_o}),
    .d({_al_u5520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] }),
    .f({_al_u5629_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Snihu6 }));
  // ../RTL/cortexm0ds_logic.v(20098)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D@C))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(B*~A*~(D@C))"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000000000100),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0100000000000100),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5632|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6_reg  (
    .a({_al_u5618_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[3]_i1[3]_o_lutinv }),
    .b({_al_u5625_o,_al_u5616_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[27]_i1[27]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqihu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[21]_i1[21]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 }),
    .mi({open_n52094,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .f({_al_u5632_o,_al_u5618_o}),
    .q({open_n52110,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 }));  // ../RTL/cortexm0ds_logic.v(20098)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(~D*A))"),
    //.LUT1("(B*~(C@D))"),
    .INIT_LUT0(16'b1100000001000000),
    .INIT_LUT1(16'b1100000000001100),
    .MODE("LOGIC"))
    \_al_u5633|_al_u5610  (
    .a({open_n52111,_al_u4423_o}),
    .b({_al_u5632_o,_al_u5609_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5992_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyhhu6 ,_al_u5523_o}),
    .f({_al_u5633_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyhhu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5634|_al_u2032  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J71iu6_lutinv ,_al_u1917_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wbkhu6 ,_al_u2032_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(C*~B*~(~D*~A))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0011000000100000),
    .MODE("LOGIC"))
    \_al_u5637|_al_u5636  (
    .a({_al_u5518_o,_al_u5523_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq0/xor_i0[1]_i1[1]_o_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 }),
    .c({_al_u5635_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 }),
    .d({_al_u5636_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u5637_o,_al_u5636_o}));
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u563|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b7  (
    .a({_al_u456_o,open_n52180}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/i_paddr [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] }),
    .mi({open_n52191,\u_cmsdk_mcu/HADDR [9]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ,_al_u462_o}),
    .q({open_n52195,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5648|_al_u5279  (
    .b({_al_u5647_o,open_n52198}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .f({_al_u5648_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2qiu6 }));
  // ../RTL/cortexm0ds_logic.v(18309)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5650|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,open_n52223}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eagax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv }),
    .mi({open_n52227,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5650_o,_al_u5812_o}),
    .q({open_n52242,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xaeax6 }));  // ../RTL/cortexm0ds_logic.v(18309)
  // ../RTL/cortexm0ds_logic.v(18217)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5651|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 ,open_n52243}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n52244}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oe7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ve7iu6 }),
    .mi({open_n52248,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5651_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oe7iu6 }),
    .q({open_n52263,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 }));  // ../RTL/cortexm0ds_logic.v(18217)
  // ../RTL/cortexm0ds_logic.v(18265)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5653|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,open_n52264}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 ,_al_u4096_o}),
    .mi({open_n52268,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktwiu6 ,_al_u5736_o}),
    .q({open_n52283,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljcax6 }));  // ../RTL/cortexm0ds_logic.v(18265)
  // ../RTL/cortexm0ds_logic.v(18331)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5654|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6_reg  (
    .a({_al_u5650_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({_al_u5651_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .c({_al_u5652_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D1aax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ktwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 }),
    .mi({open_n52294,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5654_o,_al_u5652_o}),
    .q({open_n52298,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q6fax6 }));  // ../RTL/cortexm0ds_logic.v(18331)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5657|_al_u5665  (
    .a({_al_u5649_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .b({_al_u5654_o,_al_u5657_o}),
    .c({_al_u5655_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 }),
    .d({_al_u5656_o,_al_u5664_o}),
    .f({_al_u5657_o,_al_u5665_o}));
  // ../RTL/cortexm0ds_logic.v(17806)
  EG_PHY_MSLICE #(
    //.LUT0("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101111110001000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5658|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6_reg  (
    .a({open_n52319,\u_cmsdk_mcu/HWDATA [0]}),
    .b({_al_u5260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5658_o,open_n52333}),
    .q({open_n52337,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 }));  // ../RTL/cortexm0ds_logic.v(17806)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*~B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"))
    \_al_u565|_al_u690  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n0 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5662|_al_u5660  (
    .a({open_n52360,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .b({_al_u5660_o,_al_u5067_o}),
    .c({_al_u5661_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] }),
    .d({_al_u5659_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 ,_al_u5660_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~B*~A)"),
    //.LUT1("(D*~C*B*A)"),
    .INIT_LUT0(16'b0000000000010000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"))
    \_al_u5664|_al_u5649  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaqiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K0qiu6_lutinv }),
    .b({_al_u5663_o,_al_u5291_o}),
    .c({_al_u5274_o,_al_u5648_o}),
    .d({_al_u5340_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q3qiu6 }),
    .f({_al_u5664_o,_al_u5649_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C*~(D*~B)))"),
    //.LUT1("(~B*~A*~(D*C))"),
    .INIT_LUT0(16'b0010101000001010),
    .INIT_LUT1(16'b0000000100010001),
    .MODE("LOGIC"))
    \_al_u5667|_al_u5666  (
    .a({_al_u5666_o,_al_u5020_o}),
    .b({_al_u5049_o,_al_u4865_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5665_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5667_o,_al_u5666_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5668|_al_u5050  (
    .b({_al_u5103_o,open_n52423}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 }),
    .d({_al_u5667_o,_al_u5049_o}),
    .f({_al_u5668_o,_al_u5050_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u566|_al_u567  (
    .b({open_n52450,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,_al_u566_o}),
    .f({_al_u566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b6_sel_is_13_o }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(~C*~B*~(D*A))"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(~C*~B*~(D*A))"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000000100000011),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b0000000100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5670|_al_u5672  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 ,_al_u5670_o}),
    .b({_al_u5291_o,_al_u5671_o}),
    .c({_al_u5271_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] }),
    .f({_al_u5670_o,_al_u5672_o}));
  // ../RTL/cortexm0ds_logic.v(18325)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5671|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ,open_n52499}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,open_n52500}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5671_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .q({open_n52521,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 }));  // ../RTL/cortexm0ds_logic.v(18325)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5674|_al_u5673  (
    .a({open_n52522,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 }),
    .d({_al_u5673_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtxax6 }),
    .f({_al_u5674_o,_al_u5673_o}));
  // ../RTL/cortexm0ds_logic.v(18259)
  EG_PHY_LSLICE #(
    //.LUTF0("((D@B)*(C@A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("((D@B)*(C@A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001001001000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001001001000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5676|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 ,_al_u4071_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ,_al_u4231_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxbax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 }),
    .mi({open_n52550,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .f({_al_u5676_o,_al_u5752_o}),
    .q({open_n52566,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tfcax6 }));  // ../RTL/cortexm0ds_logic.v(18259)
  // ../RTL/cortexm0ds_logic.v(18173)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5677|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6_reg  (
    .a({_al_u5672_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 }),
    .b({_al_u5674_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({_al_u5675_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5676_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vibax6 }),
    .mi({open_n52570,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .f({_al_u5677_o,_al_u5675_o}),
    .q({open_n52586,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt9ax6 }));  // ../RTL/cortexm0ds_logic.v(18173)
  // ../RTL/cortexm0ds_logic.v(20124)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000011111000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0111000011111000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5678|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/HWDATA [4]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5678_o,open_n52604}),
    .q({open_n52608,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 }));  // ../RTL/cortexm0ds_logic.v(20124)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5679|_al_u5681  (
    .a({open_n52609,_al_u5679_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ,_al_u5680_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .d({_al_u5678_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 }),
    .f({_al_u5679_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 }));
  // ../RTL/cortexm0ds_logic.v(20126)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5680|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,open_n52630}),
    .b({_al_u5067_o,open_n52631}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ,_al_u2480_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 ,\u_cmsdk_mcu/HWDATA [4]}),
    .mi({open_n52635,\u_cmsdk_mcu/HWDATA [4]}),
    .f({_al_u5680_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n152 }),
    .q({open_n52651,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Imhbx6 }));  // ../RTL/cortexm0ds_logic.v(20126)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(D*~C)))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0010101000100010),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5682|_al_u5683  (
    .a({open_n52652,_al_u5020_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0riu6 ,_al_u5682_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 ,_al_u4663_o}),
    .d({_al_u5677_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5682_o,_al_u5683_o}));
  // ../RTL/cortexm0ds_logic.v(18024)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5684|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u5683_o,_al_u1683_o}),
    .f({_al_u5684_o,open_n52689}),
    .q({open_n52693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 }));  // ../RTL/cortexm0ds_logic.v(18024)
  // ../RTL/cortexm0ds_logic.v(18023)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5685|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6_reg  (
    .b({_al_u5053_o,_al_u5103_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 }),
    .clk(XTAL1_wire),
    .d({_al_u5684_o,_al_u5685_o}),
    .f({_al_u5685_o,open_n52710}),
    .q({open_n52714,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V53qw6 }));  // ../RTL/cortexm0ds_logic.v(18023)
  // ../RTL/cortexm0ds_logic.v(19155)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110001000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1101111110001000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5687|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6_reg  (
    .a({open_n52715,\u_cmsdk_mcu/HWDATA [1]}),
    .b({_al_u5260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5687_o,open_n52733}),
    .q({open_n52737,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 }));  // ../RTL/cortexm0ds_logic.v(19155)
  // ../RTL/cortexm0ds_logic.v(17600)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5688|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6_reg  (
    .a({_al_u405_o,open_n52738}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [1]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ,_al_u2357_o}),
    .f({_al_u5688_o,open_n52753}),
    .q({open_n52757,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 }));  // ../RTL/cortexm0ds_logic.v(17600)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5691|_al_u5689  (
    .a({_al_u5689_o,_al_u5687_o}),
    .b({_al_u5690_o,_al_u5688_o}),
    .c({_al_u5067_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 ,_al_u5689_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5693|_al_u5692  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv }),
    .b({_al_u5692_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 }),
    .f({_al_u5693_o,_al_u5692_o}));
  // ../RTL/cortexm0ds_logic.v(18243)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D*~(B*A)))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~C*~(D*~(B*A)))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011111110000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111011111110000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5694|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 ,_al_u1257_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xwaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5694_o,open_n52819}),
    .q({open_n52823,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xnbax6 }));  // ../RTL/cortexm0ds_logic.v(18243)
  EG_PHY_LSLICE #(
    //.LUTF0("(A@(D*~(~C*~B)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(A@(D*~(~C*~B)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0101011010101010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0101011010101010),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5695|_al_u5402  (
    .a({open_n52824,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chkhu6 }),
    .b({open_n52825,_al_u1888_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 ,_al_u5399_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz9ax6 }),
    .f({_al_u5695_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/eq1/xor_i0[1]_i1[1]_o_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~(~B*A)))"),
    //.LUT1("(C*~B*~(D*A))"),
    .INIT_LUT0(16'b1111001000000000),
    .INIT_LUT1(16'b0001000000110000),
    .MODE("LOGIC"))
    \_al_u5697|_al_u6667  (
    .a({_al_u927_o,_al_u927_o}),
    .b({_al_u5695_o,_al_u1299_o}),
    .c({_al_u5696_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 }),
    .d({_al_u1385_o,_al_u1385_o}),
    .f({_al_u5697_o,_al_u6667_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5698|_al_u5530  (
    .a({_al_u5694_o,open_n52870}),
    .b({_al_u5697_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdbax6 ,_al_u5519_o}),
    .f({_al_u5698_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n5995_lutinv }));
  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u569|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b6  (
    .a({_al_u473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [6]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b6_sel_is_13_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b6/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .mi({open_n52894,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u569_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux3_b6/B1_0 }),
    .q({open_n52909,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [6]}));  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(C*~(D*~B)))"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(A*~(C*~(D*~B)))"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0010101000001010),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b0010101000001010),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5701|_al_u5700  (
    .a({_al_u5700_o,_al_u5020_o}),
    .b({_al_u5050_o,_al_u4581_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u5699_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9bbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u5701_o,_al_u5700_o}));
  // ../RTL/cortexm0ds_logic.v(18041)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5702|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6_reg  (
    .b({_al_u5053_o,_al_u5834_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5701_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .f({_al_u5702_o,open_n52954}),
    .q({open_n52958,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 }));  // ../RTL/cortexm0ds_logic.v(18041)
  // ../RTL/cortexm0ds_logic.v(18004)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u5705|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L18iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }),
    .c({_al_u5704_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4bax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fd7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u3885_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .mi({open_n52964,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5705_o,_al_u5704_o}),
    .q({open_n52979,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gr2qw6 }));  // ../RTL/cortexm0ds_logic.v(18004)
  // ../RTL/cortexm0ds_logic.v(19967)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(~D*~A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100101010),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5707|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6_reg  (
    .a({_al_u4035_o,_al_u4101_o}),
    .b({_al_u4101_o,_al_u4136_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 }),
    .mi({open_n52990,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .f({_al_u5707_o,_al_u5722_o}),
    .q({open_n52995,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2dbx6 }));  // ../RTL/cortexm0ds_logic.v(19967)
  // ../RTL/cortexm0ds_logic.v(19938)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~(D*B)*~(~C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0011001011111010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5709|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6_reg  (
    .a({_al_u4061_o,_al_u922_o}),
    .b({_al_u4225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ,_al_u925_o}),
    .mi({open_n53006,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .f({_al_u5709_o,_al_u926_o}),
    .q({open_n53011,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 }));  // ../RTL/cortexm0ds_logic.v(19938)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*A*(D@C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*A*(D@C))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000100010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5710|_al_u6799  (
    .a({_al_u5708_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u5709_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .c({_al_u4091_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K5hbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 }),
    .f({_al_u5710_o,_al_u6799_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(C@B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*(C@B))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0011110000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0011110000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5714|_al_u5708  (
    .a({_al_u5710_o,open_n53036}),
    .b({_al_u5711_o,_al_u4191_o}),
    .c({_al_u5712_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Apcax6 }),
    .d({_al_u5713_o,_al_u5707_o}),
    .f({_al_u5714_o,_al_u5708_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("((C@B)*(D@A))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5715|_al_u4918  (
    .a({_al_u4081_o,open_n53061}),
    .b({_al_u4131_o,_al_u4076_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 ,_al_u4081_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdebx6 ,_al_u4071_o}),
    .f({_al_u5715_o,_al_u4918_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(B*A*(D@C))"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(B*A*(D@C))"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b0000100010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5717|_al_u5576  (
    .a({_al_u5715_o,open_n53086}),
    .b({_al_u5716_o,_al_u5575_o}),
    .c({_al_u4111_o,_al_u5523_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4dax6 ,_al_u4111_o}),
    .f({_al_u5717_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9ihu6 }));
  // ../RTL/cortexm0ds_logic.v(18273)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(B*A*(D@C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0000100010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5720|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6_reg  (
    .a({_al_u5718_o,_al_u1882_o}),
    .b({_al_u5719_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .c({_al_u4056_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n53121,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .f({_al_u5720_o,_al_u2290_o}),
    .q({open_n53126,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 }));  // ../RTL/cortexm0ds_logic.v(18273)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*A*(D@B))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*A*(D@B))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0010000010000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010000010000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5721|_al_u5730  (
    .a({open_n53127,_al_u5721_o}),
    .b({_al_u5717_o,_al_u4423_o}),
    .c({_al_u5720_o,_al_u5729_o}),
    .d({_al_u5714_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlcax6 }),
    .f({_al_u5721_o,_al_u5730_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("((D@B)*(C@A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("((D@B)*(C@A))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0001001001001000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0001001001001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5726|_al_u4551  (
    .a({_al_u4116_o,open_n53152}),
    .b({_al_u4184_o,_al_u4184_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F59bx6 ,_al_u4191_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqcax6 ,_al_u4096_o}),
    .f({_al_u5726_o,_al_u4551_o}));
  // ../RTL/cortexm0ds_logic.v(18280)
  EG_PHY_LSLICE #(
    //.LUTF0("((D@B)*(C@A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("((D@B)*(C@A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001001001000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001001001000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5727|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6_reg  (
    .a({_al_u5723_o,_al_u4086_o}),
    .b({_al_u5724_o,_al_u4219_o}),
    .c({_al_u5725_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etfbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5726_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 }),
    .mi({open_n53180,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 }),
    .f({_al_u5727_o,_al_u5724_o}),
    .q({open_n53196,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q9dax6 }));  // ../RTL/cortexm0ds_logic.v(18280)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(B*A*(D@C))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000100010000000),
    .MODE("LOGIC"))
    \_al_u5729|_al_u1956  (
    .a({_al_u5727_o,open_n53197}),
    .b({_al_u5728_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfqow6 }),
    .c({_al_u4121_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Asupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U7dax6 ,_al_u1955_o}),
    .f({_al_u5729_o,_al_u1956_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*~C*B*A)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"))
    \_al_u572|_al_u571  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ,open_n53218}),
    .b({_al_u571_o,open_n53219}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .f({_al_u572_o,_al_u571_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(~D*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0011111100101010),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5731|_al_u5747  (
    .a({open_n53240,_al_u4035_o}),
    .b({open_n53241,_al_u4106_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Facax6 }),
    .d({_al_u4106_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 }),
    .f({_al_u5731_o,_al_u5747_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*(D@C))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000100010000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5732|_al_u5733  (
    .a({open_n53262,_al_u5731_o}),
    .b({open_n53263,_al_u5732_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ,_al_u4191_o}),
    .d({_al_u4126_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htbax6 }),
    .f({_al_u5732_o,_al_u5733_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(~D*~B)*~(~C*~A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(~D*~B)*~(~C*~A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111101011001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111101011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5734|_al_u5746  (
    .a({_al_u4081_o,_al_u4081_o}),
    .b({_al_u4126_o,_al_u4101_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8ebx6 }),
    .f({_al_u5734_o,_al_u5746_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*(C@A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0101101001001000),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u5735|_al_u5794  (
    .a({_al_u5733_o,_al_u4081_o}),
    .b({_al_u5734_o,_al_u4131_o}),
    .c({_al_u4035_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Daebx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 }),
    .f({_al_u5735_o,_al_u5794_o}));
  // ../RTL/cortexm0ds_logic.v(18252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(~D*~A))"),
    //.LUTF1("(~(C*B)*~(~D*~A))"),
    //.LUTG0("(~(C*B)*~(~D*~A))"),
    //.LUTG1("(~(C*B)*~(~D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100101010),
    .INIT_LUTF1(16'b0011111100101010),
    .INIT_LUTG0(16'b0011111100101010),
    .INIT_LUTG1(16'b0011111100101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5738|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6_reg  (
    .a({_al_u4136_o,_al_u4066_o}),
    .b({_al_u4225_o,_al_u4136_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 }),
    .mi({open_n53331,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .f({_al_u5738_o,_al_u5741_o}),
    .q({open_n53347,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cax6 }));  // ../RTL/cortexm0ds_logic.v(18252)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*(D@C))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(B*A*(D@C))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000100010000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5742|_al_u5771  (
    .a({_al_u5738_o,_al_u5769_o}),
    .b({_al_u5739_o,_al_u5770_o}),
    .c({_al_u5740_o,_al_u4136_o}),
    .d({_al_u5741_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 }),
    .f({_al_u5742_o,_al_u5771_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(~D*~A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1111110010101000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5745|_al_u5743  (
    .a({_al_u5737_o,_al_u4096_o}),
    .b({_al_u5742_o,_al_u4111_o}),
    .c({_al_u5743_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 }),
    .d({_al_u5744_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdcbx6 }),
    .f({_al_u5745_o,_al_u5743_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(~(C*B)*~(~D*~A))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0011111100101010),
    .MODE("LOGIC"))
    \_al_u5748|_al_u5240  (
    .a({_al_u4091_o,_al_u5238_o}),
    .b({_al_u4237_o,_al_u5239_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 }),
    .f({_al_u5748_o,_al_u5240_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~C*~B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0101010011111100),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0101010011111100),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5750|_al_u5749  (
    .a({_al_u5746_o,_al_u4091_o}),
    .b({_al_u5747_o,_al_u4101_o}),
    .c({_al_u5748_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxcbx6 }),
    .d({_al_u5749_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 }),
    .f({_al_u5750_o,_al_u5749_o}));
  // ../RTL/cortexm0ds_logic.v(19979)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5751|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6_reg  (
    .a({_al_u4076_o,open_n53436}),
    .b({_al_u4184_o,open_n53437}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5751_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .q({open_n53458,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 }));  // ../RTL/cortexm0ds_logic.v(19979)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5755|_al_u3383  (
    .a({_al_u5751_o,open_n53459}),
    .b({_al_u5752_o,open_n53460}),
    .c({_al_u5753_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7zhu6 }),
    .d({_al_u5754_o,_al_u2293_o}),
    .f({_al_u5755_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbyhu6 }));
  // ../RTL/cortexm0ds_logic.v(18245)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5756|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6_reg  (
    .a({_al_u5735_o,_al_u4423_o}),
    .b({_al_u5745_o,_al_u5756_o}),
    .c({_al_u5750_o,_al_u5758_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5755_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 }),
    .mi({open_n53484,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 }),
    .f({_al_u5756_o,_al_u5759_o}),
    .q({open_n53500,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Opbax6 }));  // ../RTL/cortexm0ds_logic.v(18245)
  // ../RTL/cortexm0ds_logic.v(19935)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(D*(C@B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0011110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5758|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6_reg  (
    .a({open_n53501,_al_u6664_o}),
    .b({_al_u4061_o,_al_u6665_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5757_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 }),
    .mi({open_n53512,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .f({_al_u5758_o,_al_u6666_o}),
    .q({open_n53517,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knbbx6 }));  // ../RTL/cortexm0ds_logic.v(19935)
  // ../RTL/cortexm0ds_logic.v(20101)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("((D@B)*(C@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0001001001001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5762|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6_reg  (
    .a({_al_u4061_o,_al_u2252_o}),
    .b({_al_u4091_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({open_n53528,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .f({_al_u5762_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jwxow6 }),
    .q({open_n53533,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3hbx6 }));  // ../RTL/cortexm0ds_logic.v(20101)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*A*~(C*B))"),
    //.LUTF1("(C*B*(D@A))"),
    //.LUTG0("(D*A*~(C*B))"),
    //.LUTG1("(C*B*(D@A))"),
    .INIT_LUTF0(16'b0010101000000000),
    .INIT_LUTF1(16'b0100000010000000),
    .INIT_LUTG0(16'b0010101000000000),
    .INIT_LUTG1(16'b0100000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5763|_al_u5723  (
    .a({_al_u4423_o,_al_u5722_o}),
    .b({_al_u5761_o,_al_u4061_o}),
    .c({_al_u5762_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Btbbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efdax6 }),
    .f({_al_u5763_o,_al_u5723_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*~(D*B))"),
    //.LUT1("(~(~D*~B)*~(C*A))"),
    .INIT_LUT0(16'b0010000010100000),
    .INIT_LUT1(16'b0101111101001100),
    .MODE("LOGIC"))
    \_al_u5765|_al_u6755  (
    .a({_al_u4081_o,_al_u6753_o}),
    .b({_al_u4191_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ,_al_u6754_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 }),
    .f({_al_u5765_o,_al_u6755_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(B*A*(D@C))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(B*A*(D@C))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000100010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5766|_al_u5333  (
    .a({_al_u5764_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u5765_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 }),
    .c({_al_u4225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 }),
    .f({_al_u5766_o,_al_u5333_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(~D*~B)*~(C*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0101111101001100),
    .MODE("LOGIC"))
    \_al_u5769|_al_u5069  (
    .a({_al_u4197_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u4231_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 }),
    .f({_al_u5769_o,_al_u5069_o}));
  // ../RTL/cmsdk_apb_uart.v(501)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u576|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2_reg  (
    .a({open_n53622,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]}),
    .b({_al_u575_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .clk(XTAL1_wire),
    .d({_al_u574_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .mi({open_n53633,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u576_o,_al_u575_o}),
    .q({open_n53637,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2 }));  // ../RTL/cmsdk_apb_uart.v(501)
  // ../RTL/cortexm0ds_logic.v(20187)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("((D@B)*(C@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001001001001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5772|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6_reg  (
    .a({_al_u4126_o,open_n53638}),
    .b({_al_u4237_o,open_n53639}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 }),
    .q({open_n53656,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 }));  // ../RTL/cortexm0ds_logic.v(20187)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5775|_al_u5773  (
    .a({_al_u5771_o,_al_u4184_o}),
    .b({_al_u5772_o,_al_u4231_o}),
    .c({_al_u5773_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7eax6 }),
    .d({_al_u5774_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 }),
    .f({_al_u5775_o,_al_u5773_o}));
  // ../RTL/cortexm0ds_logic.v(19894)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010000101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5777|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6_reg  (
    .a({_al_u4086_o,open_n53681}),
    .b({_al_u4131_o,open_n53682}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hrfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .mi({open_n53693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .f({_al_u5777_o,_al_u2129_o}),
    .q({open_n53698,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 }));  // ../RTL/cortexm0ds_logic.v(19894)
  // ../RTL/cortexm0ds_logic.v(18295)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTF1("((D@B)*(C@A))"),
    //.LUTG0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG1("((D@B)*(C@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010111000111111),
    .INIT_LUTF1(16'b0001001001001000),
    .INIT_LUTG0(16'b0010111000111111),
    .INIT_LUTG1(16'b0001001001001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5778|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6_reg  (
    .a({_al_u4056_o,_al_u4500_o}),
    .b({_al_u4116_o,_al_u4501_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J39bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9ypw6 }),
    .mi({open_n53702,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .f({_al_u5778_o,_al_u4909_o}),
    .q({open_n53718,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsdax6 }));  // ../RTL/cortexm0ds_logic.v(18295)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5780|_al_u5781  (
    .a({_al_u5776_o,_al_u5763_o}),
    .b({_al_u5777_o,_al_u5768_o}),
    .c({_al_u5778_o,_al_u5775_o}),
    .d({_al_u5779_o,_al_u5780_o}),
    .f({_al_u5780_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhhu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*(C@B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*(C@B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011110000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5784|_al_u5783  (
    .a({open_n53739,_al_u4101_o}),
    .b({_al_u4056_o,_al_u4225_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 }),
    .d({_al_u5783_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 }),
    .f({_al_u5784_o,_al_u5783_o}));
  // ../RTL/cortexm0ds_logic.v(18318)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~D*~B)*~(~C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111101011001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5785|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6_reg  (
    .a({_al_u4071_o,open_n53764}),
    .b({_al_u4136_o,open_n53765}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5785_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .q({open_n53782,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 }));  // ../RTL/cortexm0ds_logic.v(18318)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*~(~C*~A))"),
    //.LUT1("(B*A*(D@C))"),
    .INIT_LUT0(16'b1111101011001000),
    .INIT_LUT1(16'b0000100010000000),
    .MODE("LOGIC"))
    \_al_u5786|_al_u5716  (
    .a({_al_u5784_o,_al_u4035_o}),
    .b({_al_u5785_o,_al_u4237_o}),
    .c({_al_u4237_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B9jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 }),
    .f({_al_u5786_o,_al_u5716_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(C@B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*(C@B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0011110000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0011110000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5787|_al_u5737  (
    .b({open_n53805,_al_u4197_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hjgax6 }),
    .d({_al_u4096_o,_al_u5736_o}),
    .f({_al_u5787_o,_al_u5737_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5791|_al_u5790  (
    .a({_al_u5786_o,_al_u4035_o}),
    .b({_al_u5788_o,_al_u4121_o}),
    .c({_al_u5789_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 }),
    .d({_al_u5790_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 }),
    .f({_al_u5791_o,_al_u5790_o}));
  // ../RTL/cortexm0ds_logic.v(18319)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(~D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111100101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5792|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6_reg  (
    .a({_al_u4101_o,open_n53854}),
    .b({_al_u4126_o,open_n53855}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fj8ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zycbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u5792_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .q({open_n53872,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 }));  // ../RTL/cortexm0ds_logic.v(18319)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5797|_al_u5796  (
    .a({open_n53873,_al_u4131_o}),
    .b({_al_u5795_o,_al_u4136_o}),
    .c({_al_u5796_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 }),
    .d({_al_u5794_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 }),
    .f({_al_u5797_o,_al_u5796_o}));
  // ../RTL/cortexm0ds_logic.v(18322)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(C@B))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011110000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5800|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6_reg  (
    .a({_al_u5793_o,open_n53898}),
    .b({_al_u5797_o,_al_u4106_o}),
    .c({_al_u5798_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5799_o,_al_u5792_o}),
    .mi({open_n53909,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .f({_al_u5800_o,_al_u5793_o}),
    .q({open_n53914,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxeax6 }));  // ../RTL/cortexm0ds_logic.v(18322)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("((D@B)*(C@A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("((D@B)*(C@A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001001001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001001001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5805|_al_u5317  (
    .a({_al_u4219_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u4231_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1fax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y2fax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 }),
    .f({_al_u5805_o,_al_u5317_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5806|_al_u6798  (
    .a({_al_u5802_o,open_n53939}),
    .b({_al_u5803_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u5804_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztgbx6 }),
    .d({_al_u5805_o,_al_u6797_o}),
    .f({_al_u5806_o,_al_u6798_o}));
  // ../RTL/cortexm0ds_logic.v(18312)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*A*~(D*C))"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000100010),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5809|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6_reg  (
    .a({open_n53964,_al_u5760_o}),
    .b({open_n53965,_al_u5782_o}),
    .c({_al_u5808_o,_al_u5809_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5801_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 }),
    .mi({open_n53976,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .f({_al_u5809_o,_al_u5810_o}),
    .q({open_n53981,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Peeax6 }));  // ../RTL/cortexm0ds_logic.v(18312)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u581|_al_u4565  (
    .a({open_n53982,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]}),
    .d({_al_u580_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}),
    .f({_al_u581_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n12_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(D*~(C*~B*A))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"))
    \_al_u5839|_al_u5838  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiaju6 ,_al_u696_o}),
    .b({_al_u4351_o,_al_u932_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejaju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejaju6_lutinv }));
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u583|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b6  (
    .a({open_n54027,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .b({open_n54028,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}),
    .c({_al_u582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5]}),
    .clk(XTAL1_wire),
    .d({_al_u581_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}),
    .mi({open_n54033,\u_cmsdk_mcu/HADDR [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ,_al_u582_o}),
    .q({open_n54048,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_MSLICE #(
    //.LUT0("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100100011111000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5841|_al_u5840  (
    .a({open_n54049,_al_u1344_o}),
    .b({open_n54050,_al_u2403_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ,_al_u3826_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5842|_al_u929  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nkaju6_lutinv ,open_n54073}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUTF1("(A*~(~B*~(~D*C)))"),
    //.LUTG0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUTG1("(A*~(~B*~(~D*C)))"),
    .INIT_LUTF0(16'b0111111101001100),
    .INIT_LUTF1(16'b1000100010101000),
    .INIT_LUTG0(16'b0111111101001100),
    .INIT_LUTG1(16'b1000100010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5845|_al_u5843  (
    .a({_al_u5843_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({_al_u5845_o,_al_u5843_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~C*~B*D)"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"))
    \_al_u5847|_al_u5846  (
    .a({open_n54118,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 }));
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    //.LUT1("(~D*~(~B*~(~C*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110010001000100),
    .INIT_LUT1(16'b0000000011001101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u584|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hz0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qc3pw6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u584_o,\u_cmsdk_mcu/HADDR [1]}),
    .q({open_n54155,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [1]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*A))"),
    //.LUT1("(D*~(B*~(~C*~A)))"),
    .INIT_LUT0(16'b0100110001011111),
    .INIT_LUT1(16'b0011011100000000),
    .MODE("LOGIC"))
    \_al_u5852|_al_u5851  (
    .a({_al_u5850_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Difiu6 }),
    .b({_al_u5851_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u5851_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*~B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0100000001010000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5853|_al_u5855  (
    .a({open_n54176,_al_u5845_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u2281_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32],_al_u5853_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N45ju6 ,_al_u5854_o}),
    .f({_al_u5853_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5858|_al_u5857  (
    .a({open_n54197,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u5848_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31],n1[12]}),
    .d({_al_u5857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] }),
    .f({_al_u5858_o,_al_u5857_o}));
  // ../RTL/cmsdk_ahb_to_iop.v(69)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(D*C*B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u585|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_ahb_to_gpio/IOSEL_reg  (
    .a({_al_u584_o,open_n54222}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ,open_n54223}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio1_hsel }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u585_o,open_n54237}),
    .q({open_n54241,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL }));  // ../RTL/cmsdk_ahb_to_iop.v(69)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))"),
    //.LUTF1("(B*~(~D*C*~A))"),
    //.LUTG0("(A*~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))"),
    //.LUTG1("(B*~(~D*C*~A))"),
    .INIT_LUTF0(16'b0010101000001000),
    .INIT_LUTF1(16'b1100110010001100),
    .INIT_LUTG0(16'b0010101000001000),
    .INIT_LUTG1(16'b1100110010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5860|_al_u5856  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30]}),
    .b({_al_u5859_o,_al_u1541_o}),
    .c({_al_u1541_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({_al_u5860_o,_al_u5856_o}));
  // ../RTL/cortexm0ds_logic.v(17906)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~C*B*~A)"),
    //.LUTF1("(~D*C*~B*A)"),
    //.LUTG0("~(D*~C*B*~A)"),
    //.LUTG1("(~D*C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101111111111),
    .INIT_LUTF1(16'b0000000000100000),
    .INIT_LUTG0(16'b1111101111111111),
    .INIT_LUTG1(16'b0000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5861|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ykzpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 ,_al_u7092_o}),
    .b({_al_u5856_o,_al_u7117_o}),
    .c({_al_u5860_o,_al_u5856_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ,_al_u5860_o}),
    .f({_al_u5861_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .q({open_n54286,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[28] }));  // ../RTL/cortexm0ds_logic.v(17906)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1100100011000000),
    .MODE("LOGIC"))
    \_al_u5862|_al_u1534  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29],open_n54287}),
    .b({_al_u1533_o,open_n54288}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ,_al_u1348_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ,_al_u1533_o}),
    .f({_al_u5862_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [29]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000000100000011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5864|_al_u5863  (
    .a({open_n54309,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u5848_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30],n1[11]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J77ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] }),
    .f({_al_u5864_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J77ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*(C@B)))"),
    //.LUT1("(C*~A*~(D*~B))"),
    .INIT_LUT0(16'b1000001010101010),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"))
    \_al_u5865|_al_u5866  (
    .a({_al_u5862_o,_al_u5865_o}),
    .b({_al_u2429_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29]}),
    .c({_al_u5864_o,_al_u1533_o}),
    .d({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({_al_u5865_o,_al_u5866_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5869|_al_u5868  (
    .a({open_n54350,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5868_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[7]}),
    .d({_al_u2261_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26]}),
    .f({_al_u5869_o,_al_u5868_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(D*~C)))"),
    //.LUT1("(B*~(~A*~(D*~C)))"),
    .INIT_LUT0(16'b1000110010001000),
    .INIT_LUT1(16'b1000110010001000),
    .MODE("LOGIC"))
    \_al_u586|_al_u592  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv }),
    .b({_al_u585_o,_al_u591_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n39 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5871|_al_u5867  (
    .a({open_n54395,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25]}),
    .b({open_n54396,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mi8ju6_lutinv }),
    .c({_al_u5870_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yh8ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5871_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yh8ju6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u5875|_al_u5874  (
    .a({open_n54421,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 }),
    .b({_al_u5848_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .d({_al_u5874_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o }),
    .f({_al_u5875_o,_al_u5874_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5877|_al_u5876  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .d({_al_u5875_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wy4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5878|_al_u5977  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wy4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pa7ju6 }),
    .f({_al_u5878_o,_al_u5977_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~A*~(D*~C))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b0100000001000100),
    .MODE("LOGIC"))
    \_al_u5879|_al_u5873  (
    .a({_al_u5873_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0]}),
    .b({_al_u5878_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv }),
    .c({_al_u1882_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .d({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv }),
    .f({_al_u5879_o,_al_u5873_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(~D*~(~B*~(~C*A)))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(~D*~(~B*~(~C*A)))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0000000011001110),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0000000011001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u587|_al_u4550  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [0],open_n54506}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [1],_al_u4549_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSIZE [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .f({_al_u587_o,_al_u4550_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(~C*~(D*~A)))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(~C*~(D*~A)))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1100010011000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1100010011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5880|_al_u5844  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0],open_n54531}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Go0iu6_lutinv ,open_n54532}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 }),
    .f({_al_u5880_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(18973)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5881|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1yax6_reg  (
    .c({_al_u5880_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5879_o,_al_u7028_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .q({open_n54577,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] }));  // ../RTL/cortexm0ds_logic.v(18973)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5884|_al_u5883  (
    .a({open_n54578,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5883_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_9 }),
    .f({_al_u5884_o,_al_u5883_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C@(A*~(D*~B)))"),
    //.LUTF1("(B*~(D*C*A))"),
    //.LUTG0("~(C@(A*~(D*~B)))"),
    //.LUTG1("(B*~(D*C*A))"),
    .INIT_LUTF0(16'b1000011110100101),
    .INIT_LUTF1(16'b0100110011001100),
    .INIT_LUTG0(16'b1000011110100101),
    .INIT_LUTG1(16'b0100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5885|_al_u2465  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ,_al_u2464_o}),
    .b({_al_u5884_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I28ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv ,_al_u2398_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ,_al_u2412_o}),
    .f({_al_u5885_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5886|_al_u5882  (
    .a({open_n54627,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 }),
    .b({open_n54628,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N18ju6_lutinv }),
    .c({_al_u5885_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z08ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5886_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z08ju6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(18764)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5887|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wrmax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ibliu6 ,_al_u6989_o}),
    .c({_al_u5886_o,_al_u5886_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5872_o,_al_u6969_o}),
    .f({_al_u5887_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .q({open_n54671,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[9] }));  // ../RTL/cortexm0ds_logic.v(18764)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(D*C*B*~A)"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b0100000000000000),
    .MODE("LOGIC"))
    \_al_u588|_al_u593  (
    .a({_al_u587_o,_al_u587_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/IOSEL ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE }),
    .f({_al_u588_o,_al_u593_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u5890|_al_u5889  (
    .a({open_n54692,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5889_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7]}),
    .d({_al_u1952_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_6 }),
    .f({_al_u5890_o,_al_u5889_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u5892|_al_u5888  (
    .a({open_n54713,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 }),
    .b({open_n54714,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk6ju6_lutinv }),
    .c({_al_u5891_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5888_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5892_o,_al_u5888_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUT1("(A*~(~B*~(~D*C)))"),
    .INIT_LUT0(16'b0111111101001100),
    .INIT_LUT1(16'b1000100010101000),
    .MODE("LOGIC"))
    \_al_u5894|_al_u5893  (
    .a({_al_u5893_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24],_al_u1493_o}),
    .c({_al_u1493_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({_al_u5894_o,_al_u5893_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~(D*A))"),
    //.LUT1("(C*~A*~(D*~B))"),
    .INIT_LUT0(16'b0000000100000011),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"))
    \_al_u5896|_al_u5895  (
    .a({_al_u5894_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u2439_o,_al_u5848_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ww6ju6 ,n1[6]}),
    .d({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25]}),
    .f({_al_u5896_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ww6ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*~B))"),
    //.LUT1("(B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0100000001010000),
    .INIT_LUT1(16'b1100100011000000),
    .MODE("LOGIC"))
    \_al_u5897|_al_u5900  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28],_al_u5897_o}),
    .b({_al_u1525_o,_al_u2420_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 ,_al_u5899_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tt4ju6_lutinv ,_al_u5854_o}),
    .f({_al_u5897_o,_al_u5900_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5899|_al_u5898  (
    .a({open_n54795,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u5848_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29],n1[10]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] }),
    .f({_al_u5899_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ok7ju6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u589|_al_u4566  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ,_al_u4566_o}));
  // ../RTL/cortexm0ds_logic.v(17217)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(A*~(D*(C@B)))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(A*~(D*(C@B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b1000001010101010),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b1000001010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5901|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uqipw6_reg  (
    .a({_al_u5900_o,open_n54848}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28],open_n54849}),
    .c({_al_u1525_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ,_al_u7122_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .q({open_n54870,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[28] }));  // ../RTL/cortexm0ds_logic.v(17217)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5904|_al_u5903  (
    .a({open_n54871,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5903_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[9]}),
    .d({_al_u2447_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28]}),
    .f({_al_u5904_o,_al_u5903_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u5906|_al_u5902  (
    .a({open_n54896,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27]}),
    .b({open_n54897,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F57ju6_lutinv }),
    .c({_al_u5905_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R47ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R47ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5909|_al_u5908  (
    .a({open_n54918,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5908_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[8]}),
    .d({_al_u2455_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27]}),
    .f({_al_u5909_o,_al_u5908_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u590|_al_u594  (
    .b({_al_u588_o,_al_u593_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n26_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n24_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n34 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5911|_al_u5907  (
    .a({open_n54965,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26]}),
    .b({open_n54966,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E17ju6_lutinv }),
    .c({_al_u5910_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q07ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5911_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q07ju6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17900)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5912|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8zpw6_reg  (
    .a({_al_u5896_o,open_n54991}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kgoiu6 ,open_n54992}),
    .c({_al_u5906_o,_al_u5896_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5911_o,_al_u7101_o}),
    .f({_al_u5912_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .q({open_n55013,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[22] }));  // ../RTL/cortexm0ds_logic.v(17900)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5913|_al_u5872  (
    .b({_al_u5892_o,_al_u5866_o}),
    .c({_al_u5912_o,_al_u5871_o}),
    .d({_al_u5887_o,_al_u5861_o}),
    .f({_al_u5913_o,_al_u5872_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u5916|_al_u5915  (
    .a({open_n55040,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5915_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_8 }),
    .f({_al_u5916_o,_al_u5915_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C@(A*~(D*~B)))"),
    //.LUT1("(C*~(D*~B*A))"),
    .INIT_LUT0(16'b1000011110100101),
    .INIT_LUT1(16'b1101000011110000),
    .MODE("LOGIC"))
    \_al_u5917|_al_u2879  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 ,_al_u2878_o}),
    .b({_al_u1608_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz7ju6 }),
    .c({_al_u5916_o,_al_u2398_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ,_al_u2412_o}),
    .f({_al_u5917_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100001001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100001001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5918|_al_u5914  (
    .a({open_n55081,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 }),
    .b({open_n55082,_al_u1608_o}),
    .c({_al_u5917_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs7ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5918_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs7ju6_lutinv }));
  // ../RTL/cmsdk_ahb_to_iop.v(69)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(D*C*B*~A)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(D*C*B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u591|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/IOSEL_reg  (
    .a({_al_u584_o,open_n55107}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL ,open_n55108}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOTRANS ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_hsel }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u591_o,open_n55126}),
    .q({open_n55130,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOSEL }));  // ../RTL/cmsdk_ahb_to_iop.v(69)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u5921|_al_u5920  (
    .a({open_n55131,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5920_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17]}),
    .d({_al_u2289_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_16 }),
    .f({_al_u5921_o,_al_u5920_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u5923|_al_u5919  (
    .a({open_n55152,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 }),
    .b({open_n55153,_al_u1429_o}),
    .c({_al_u5922_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5919_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 ,_al_u5919_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5926|_al_u5925  (
    .a({open_n55174,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5925_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[0]}),
    .d({_al_u2208_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19]}),
    .f({_al_u5926_o,_al_u5925_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u5928|_al_u5924  (
    .a({open_n55199,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 }),
    .b({open_n55200,_al_u1445_o}),
    .c({_al_u5927_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5924_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 ,_al_u5924_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5931|_al_u5930  (
    .a({open_n55221,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5930_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13]}),
    .d({_al_u2084_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_12 }),
    .f({_al_u5931_o,_al_u5930_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100001001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100001001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5933|_al_u5929  (
    .a({open_n55246,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 }),
    .b({open_n55247,_al_u1397_o}),
    .c({_al_u5932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5929_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5933_o,_al_u5929_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u5934|_al_u7027  (
    .a({_al_u5918_o,open_n55272}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 ,_al_u7023_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 }),
    .d({_al_u5933_o,_al_u6846_o}),
    .f({_al_u5934_o,_al_u7027_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~(D*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000100000011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u5937|_al_u5936  (
    .a({open_n55293,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5936_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[1]}),
    .d({_al_u2217_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20]}),
    .f({_al_u5937_o,_al_u5936_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100001001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100001001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5939|_al_u5935  (
    .a({open_n55314,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 }),
    .b({open_n55315,_al_u1453_o}),
    .c({_al_u5938_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5935_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 ,_al_u5935_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~(D*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000100000011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u5942|_al_u5941  (
    .a({open_n55340,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5941_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[2]}),
    .d({_al_u2225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21]}),
    .f({_al_u5942_o,_al_u5941_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u5944|_al_u5940  (
    .a({open_n55361,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 }),
    .b({open_n55362,_al_u1461_o}),
    .c({_al_u5943_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5940_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 ,_al_u5940_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5947|_al_u5946  (
    .a({open_n55383,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5946_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[3]}),
    .d({_al_u2235_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22]}),
    .f({_al_u5947_o,_al_u5946_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u5949|_al_u5945  (
    .a({open_n55408,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 }),
    .b({open_n55409,_al_u1469_o}),
    .c({_al_u5948_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5945_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 ,_al_u5945_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5952|_al_u5951  (
    .a({open_n55430,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5951_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14]}),
    .d({_al_u2106_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_13 }),
    .f({_al_u5952_o,_al_u5951_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100001001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100001001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5954|_al_u5950  (
    .a({open_n55455,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 }),
    .b({open_n55456,_al_u1405_o}),
    .c({_al_u5953_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u5950_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5954_o,_al_u5950_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5956|_al_u5955  (
    .a({open_n55481,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y4miu6 }),
    .b({_al_u5934_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1miu6 }),
    .c({_al_u5955_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 }),
    .d({_al_u5913_o,_al_u5954_o}),
    .f({_al_u5956_o,_al_u5955_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUT1("(A*~(~B*~(~D*C)))"),
    .INIT_LUT0(16'b0111111101001100),
    .INIT_LUT1(16'b1000100010101000),
    .MODE("LOGIC"))
    \_al_u5958|_al_u5957  (
    .a({_al_u5957_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3],_al_u1592_o}),
    .c({_al_u1592_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({_al_u5958_o,_al_u5957_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u5959|_al_u2793  (
    .b({_al_u5848_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlliu6 ,_al_u1299_o}),
    .f({_al_u5959_o,_al_u2793_o}));
  // ../RTL/cmsdk_apb_uart.v(377)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u595|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_tick_reg  (
    .b({open_n55546,_al_u556_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ,_al_u557_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n48 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ,_al_u555_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n48 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i }),
    .q({open_n55562,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK }));  // ../RTL/cmsdk_apb_uart.v(377)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(C@B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~D*(C@B))"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0000000000111100),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000000000111100),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5960|_al_u3243  (
    .b({_al_u5959_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9mpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqkax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ,_al_u2783_o}),
    .f({_al_u5960_o,_al_u3243_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(D*~B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(C*~A*~(D*~B))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0100000001010000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5961|_al_u5962  (
    .a({open_n55589,_al_u5958_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u1925_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4],_al_u5961_o}),
    .d({_al_u5960_o,_al_u5854_o}),
    .f({_al_u5961_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUTF1("(A*~(~B*~(~D*C)))"),
    //.LUTG0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUTG1("(A*~(~B*~(~D*C)))"),
    .INIT_LUTF0(16'b0111111101001100),
    .INIT_LUTF1(16'b1000100010101000),
    .INIT_LUTG0(16'b0111111101001100),
    .INIT_LUTG1(16'b1000100010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5964|_al_u5963  (
    .a({_al_u5963_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5],_al_u1600_o}),
    .c({_al_u1600_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({_al_u5964_o,_al_u5963_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5966|_al_u5965  (
    .a({open_n55638,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u5848_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I46ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_5 }),
    .f({_al_u5966_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I46ju6 }));
  // ../RTL/cortexm0ds_logic.v(18902)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(C*~A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5967|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zduax6_reg  (
    .a({_al_u5964_o,open_n55659}),
    .b({_al_u1943_o,open_n55660}),
    .c({_al_u5966_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5854_o,_al_u7045_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .q({open_n55677,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] }));  // ../RTL/cortexm0ds_logic.v(18902)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u5970|_al_u5969  (
    .a({open_n55678,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u5969_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8]}),
    .d({_al_u1961_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_7 }),
    .f({_al_u5970_o,_al_u5969_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(B*~(D*~C*A))"),
    //.LUTG0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(B*~(D*~C*A))"),
    .INIT_LUTF0(16'b0000100001001100),
    .INIT_LUTF1(16'b1100010011001100),
    .INIT_LUTG0(16'b0000100001001100),
    .INIT_LUTG1(16'b1100010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5971|_al_u5968  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 }),
    .b({_al_u5970_o,_al_u1616_o}),
    .c({_al_u1616_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u5971_o,_al_u5968_o}));
  // ../RTL/cortexm0ds_logic.v(17631)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5972|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvrpw6_reg  (
    .c({_al_u5971_o,_al_u5972_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5968_o,_al_u7053_o}),
    .f({_al_u5972_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .q({open_n55743,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[7] }));  // ../RTL/cortexm0ds_logic.v(17631)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUTF1("(A*~(~B*~(~D*C)))"),
    //.LUTG0("~(~D*~((C*A))*~(B)+~D*(C*A)*~(B)+~(~D)*(C*A)*B+~D*(C*A)*B)"),
    //.LUTG1("(A*~(~B*~(~D*C)))"),
    .INIT_LUTF0(16'b0111111101001100),
    .INIT_LUTF1(16'b1000100010101000),
    .INIT_LUTG0(16'b0111111101001100),
    .INIT_LUTG1(16'b1000100010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5974|_al_u5973  (
    .a({_al_u5973_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1],_al_u1354_o}),
    .c({_al_u1354_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .f({_al_u5974_o,_al_u5973_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~D*~B*~(C*A))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~D*~B*~(C*A))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000000010011),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5976|_al_u5975  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T05ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rb7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rskax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pa7ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rb7ju6 }));
  // ../RTL/cortexm0ds_logic.v(18752)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(C*~A*~(D*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5978|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X3max6_reg  (
    .a({_al_u5974_o,open_n55792}),
    .b({_al_u1968_o,open_n55793}),
    .c({_al_u5977_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u5854_o,_al_u7057_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .q({open_n55810,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[1] }));  // ../RTL/cortexm0ds_logic.v(18752)
  // ../RTL/cortexm0ds_logic.v(18826)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u5979|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z6qax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 ,open_n55811}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lokiu6 ,open_n55812}),
    .c({_al_u5972_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkkiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bpliu6 ,_al_u7036_o}),
    .f({_al_u5979_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .q({open_n55829,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[3] }));  // ../RTL/cortexm0ds_logic.v(18826)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b1101111011010100),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1101111011010100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5981|_al_u5980  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [2],open_n55830}),
    .b({_al_u5980_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 }),
    .c({_al_u1581_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ,_al_u1581_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am5ju6_lutinv ,_al_u5980_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~(D*A))"),
    //.LUT1("(~D*~A*~(C*B))"),
    .INIT_LUT0(16'b0000000100000011),
    .INIT_LUT1(16'b0000000000010101),
    .MODE("LOGIC"))
    \_al_u5983|_al_u5849  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk5ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I55ju6 }),
    .b({_al_u5848_o,_al_u5848_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_control_o ,n1[13]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] }),
    .f({_al_u5983_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N45ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*~(D*~B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b1000000010100000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u5985|_al_u5986  (
    .a({open_n55875,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am5ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u1916_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3],_al_u5985_o}),
    .d({_al_u5984_o,_al_u5854_o}),
    .f({_al_u5985_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5987|_al_u6210  (
    .a({open_n55896,_al_u6194_o}),
    .b({_al_u5979_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cgkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 }),
    .d({_al_u5956_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 }),
    .f({_al_u5987_o,_al_u6210_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("~(C*~D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b1111111100001111),
    .MODE("LOGIC"))
    \_al_u598|_al_u597  (
    .a({open_n55917,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 }),
    .b({open_n55918,uart0_txen_pad}),
    .c({_al_u597_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ,_al_u597_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C@B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~(C@B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011000011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011000011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5990|_al_u6006  (
    .b({open_n55941,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u5988_o,_al_u5988_o}),
    .f({_al_u5990_o,_al_u6006_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B@(C*~D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B@(C*~D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100110000111100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100110000111100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5992|_al_u5998  (
    .b({open_n55968,_al_u5991_o}),
    .c({_al_u5991_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u5990_o,_al_u5990_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ,_al_u5998_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B@(C*~D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100110000111100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5994|_al_u6039  (
    .b({open_n55995,_al_u5993_o}),
    .c({_al_u5993_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv ,_al_u6039_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B@(C*~D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B@(C*~D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100110000111100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100110000111100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5996|_al_u6038  (
    .b({open_n56018,_al_u5995_o}),
    .c({_al_u5995_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J43ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(C@B))"),
    //.LUTF1("(A*~(C@(D*~B)))"),
    //.LUTG0("(~D*(C@B))"),
    //.LUTG1("(A*~(C@(D*~B)))"),
    .INIT_LUTF0(16'b0000000000111100),
    .INIT_LUTF1(16'b0010100000001010),
    .INIT_LUTG0(16'b0000000000111100),
    .INIT_LUTG1(16'b0010100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6000|_al_u6002  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ,open_n56043}),
    .b({_al_u5988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,_al_u5988_o}),
    .f({_al_u6000_o,_al_u6002_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(C*B)))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1110101000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u6001|_al_u6947  (
    .a({open_n56068,_al_u6011_o}),
    .b({open_n56069,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 }),
    .c({_al_u6000_o,_al_u6021_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ,_al_u6817_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 ,_al_u6947_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6005|_al_u6004  (
    .a({open_n56090,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 }),
    .b({_al_u6004_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6005_o,_al_u6004_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6007|_al_u770  (
    .b({_al_u6006_o,open_n56113}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 }),
    .d({_al_u6005_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6007_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6009|_al_u6008  (
    .a({open_n56134,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 }),
    .b({_al_u6008_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6009_o,_al_u6008_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u600|_al_u564  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PWRITE ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_apb_slave_mux/n4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/apb_tran_end }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6010|_al_u6122  (
    .b({_al_u6006_o,_al_u6006_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 }),
    .d({_al_u6009_o,_al_u6121_o}),
    .f({_al_u6010_o,_al_u6122_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*C*~B))"),
    //.LUT1("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b1000101010101010),
    .INIT_LUT1(16'b0001000100000101),
    .MODE("LOGIC"))
    \_al_u6011|_al_u6003  (
    .a({_al_u6003_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lolow6 }),
    .b({_al_u6007_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .c({_al_u6010_o,_al_u5998_o}),
    .d({_al_u5998_o,_al_u6002_o}),
    .f({_al_u6011_o,_al_u6003_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b1011000100000000),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6012|_al_u5999  (
    .a({open_n56231,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kupow6_lutinv }),
    .c({_al_u5990_o,_al_u5998_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5oow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6014|_al_u6013  (
    .a({open_n56252,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 }),
    .b({_al_u6013_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6014_o,_al_u6013_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6015|_al_u866  (
    .b({_al_u6006_o,open_n56275}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 }),
    .d({_al_u6014_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6015_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6017|_al_u6016  (
    .a({open_n56296,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 }),
    .b({_al_u6016_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6017_o,_al_u6016_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6018|_al_u842  (
    .b({_al_u6006_o,open_n56323}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 }),
    .d({_al_u6017_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6018_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [6]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*A))"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(~(D*~B)*~(C*A))"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b0100110001011111),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b0100110001011111),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6021|_al_u6020  (
    .a({open_n56344,_al_u1813_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqpow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u6021_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xqpow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"))
    \_al_u6022|_al_u6019  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv ,_al_u6018_o}),
    .c({_al_u6021_o,_al_u5998_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5oow6 ,_al_u6015_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6024|_al_u6023  (
    .a({open_n56391,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 }),
    .b({_al_u6023_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6024_o,_al_u6023_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6029|_al_u6028  (
    .a({open_n56412,_al_u823_o}),
    .b({_al_u6028_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6029_o,_al_u6028_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~(B@A))"),
    //.LUTF1("(~B*~(A*~(D*~C)))"),
    //.LUTG0("(D*~C*~(B@A))"),
    //.LUTG1("(~B*~(A*~(D*~C)))"),
    .INIT_LUTF0(16'b0000100100000000),
    .INIT_LUTF1(16'b0001001100010001),
    .INIT_LUTG0(16'b0000100100000000),
    .INIT_LUTG1(16'b0001001100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6031|_al_u6027  (
    .a({_al_u6026_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .b({_al_u6027_o,_al_u5998_o}),
    .c({_al_u6030_o,_al_u6021_o}),
    .d({_al_u5998_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ,_al_u6027_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6033|_al_u6032  (
    .a({open_n56457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 }),
    .b({_al_u6032_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6033_o,_al_u6032_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6034|_al_u806  (
    .b({_al_u6002_o,open_n56484}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 }),
    .d({_al_u6033_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6034_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [25]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6035|_al_u6030  (
    .b({_al_u6034_o,_al_u6002_o}),
    .c({_al_u5998_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 }),
    .d({_al_u6030_o,_al_u6029_o}),
    .f({_al_u6035_o,_al_u6030_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~((D*A))+B*C*~((D*A))+~(B)*C*(D*A)+B*C*(D*A))"),
    //.LUT1("(D*~C*B*~A)"),
    .INIT_LUT0(16'b0001101100110011),
    .INIT_LUT1(16'b0000010000000000),
    .MODE("LOGIC"))
    \_al_u6037|_al_u6036  (
    .a({_al_u6011_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ,_al_u6035_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ,_al_u6021_o}),
    .d({_al_u6036_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u6037_o,_al_u6036_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6040|_al_u6129  (
    .b({open_n56553,_al_u6039_o}),
    .c({_al_u6039_o,_al_u6045_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv }),
    .f({_al_u6040_o,_al_u6129_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(C*~(B*D))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"))
    \_al_u6041|_al_u3572  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Svzhu6 ,_al_u932_o}),
    .c({_al_u932_o,_al_u2403_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvzhu6 ,_al_u906_o}),
    .f({_al_u6041_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rvniu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~C*~A*~(D*~B))"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000010000000101),
    .MODE("LOGIC"))
    \_al_u6044|_al_u6043  (
    .a({_al_u6041_o,_al_u607_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwzhu6 ,_al_u6042_o}),
    .c({_al_u6043_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u932_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1kpw6 }),
    .f({_al_u6044_o,_al_u6043_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6046|_al_u6100  (
    .b({open_n56618,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv }),
    .c({_al_u6045_o,_al_u6045_o}),
    .d({_al_u6040_o,_al_u6040_o}),
    .f({_al_u6046_o,_al_u6100_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6048|_al_u6131  (
    .c({_al_u6039_o,_al_u6039_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6049|_al_u6848  (
    .c({_al_u6045_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ,_al_u6049_o}),
    .f({_al_u6049_o,_al_u6848_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6051|_al_u6050  (
    .b({open_n56697,_al_u604_o}),
    .c({_al_u6050_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u6047_o,_al_u6049_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ,_al_u6050_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6053|_al_u6052  (
    .a({open_n56718,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 }),
    .b({_al_u6052_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6053_o,_al_u6052_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6054|_al_u764  (
    .b({_al_u6002_o,open_n56745}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 }),
    .d({_al_u6053_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6054_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [19]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6056|_al_u6055  (
    .a({open_n56770,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 }),
    .b({_al_u6055_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6056_o,_al_u6055_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6057|_al_u776  (
    .b({_al_u6006_o,open_n56793}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 }),
    .d({_al_u6056_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6057_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [20]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6058|_al_u6893  (
    .b({open_n56816,_al_u6054_o}),
    .c({_al_u6057_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .d({_al_u6054_o,_al_u6892_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6060|_al_u6059  (
    .a({open_n56837,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 }),
    .b({_al_u6059_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6060_o,_al_u6059_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6063|_al_u6062  (
    .a({open_n56858,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 }),
    .b({_al_u6062_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6063_o,_al_u6062_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6064|_al_u758  (
    .b({_al_u6006_o,open_n56885}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 }),
    .d({_al_u6063_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6064_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(~D*C*B*A)"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b0000000010000000),
    .MODE("LOGIC"))
    \_al_u6065|_al_u6061  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ,open_n56910}),
    .b({_al_u6061_o,_al_u6006_o}),
    .c({_al_u6064_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 }),
    .d({_al_u5998_o,_al_u6060_o}),
    .f({_al_u6065_o,_al_u6061_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6067|_al_u6066  (
    .a({open_n56931,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 }),
    .b({_al_u6066_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6067_o,_al_u6066_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6068|_al_u728  (
    .b({_al_u6006_o,open_n56958}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 }),
    .d({_al_u6067_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6068_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [13]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6070|_al_u6069  (
    .a({open_n56983,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 }),
    .b({_al_u6069_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6070_o,_al_u6069_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6072|_al_u6071  (
    .b({open_n57006,_al_u6002_o}),
    .c({_al_u6071_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 }),
    .d({_al_u6068_o,_al_u6070_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ,_al_u6071_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6074|_al_u6073  (
    .a({open_n57027,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 }),
    .b({_al_u6073_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6074_o,_al_u6073_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6075|_al_u722  (
    .b({_al_u6002_o,open_n57050}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 }),
    .d({_al_u6074_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6075_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [12]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~A*~(D*B)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~(~A*~(D*B)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1110000010100000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1110000010100000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6076|_al_u6096  (
    .a({open_n57075,_al_u6065_o}),
    .b({open_n57076,_al_u6076_o}),
    .c({_al_u6075_o,_al_u6094_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ,_al_u6095_o}),
    .f({_al_u6076_o,_al_u6096_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6078|_al_u6077  (
    .a({open_n57101,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 }),
    .b({_al_u6077_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6078_o,_al_u6077_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6079|_al_u740  (
    .b({_al_u6006_o,open_n57128}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 }),
    .d({_al_u6078_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6079_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [15]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6081|_al_u6080  (
    .a({open_n57149,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 }),
    .b({_al_u6080_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6081_o,_al_u6080_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6082|_al_u848  (
    .b({_al_u6002_o,open_n57176}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 }),
    .d({_al_u6081_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6082_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [9]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6085|_al_u6084  (
    .a({open_n57201,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 }),
    .b({_al_u6084_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6085_o,_al_u6084_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u6087|_al_u6086  (
    .b({_al_u6086_o,_al_u6006_o}),
    .c({_al_u5998_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 }),
    .d({_al_u6064_o,_al_u6085_o}),
    .f({_al_u6087_o,_al_u6086_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6089|_al_u6088  (
    .a({open_n57244,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 }),
    .b({_al_u6088_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6089_o,_al_u6088_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u608|_al_u5848  (
    .b({_al_u607_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u606_o,_al_u606_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ,_al_u5848_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6090|_al_u752  (
    .b({_al_u6006_o,open_n57289}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 }),
    .d({_al_u6089_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6092|_al_u6091  (
    .a({open_n57314,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 }),
    .b({_al_u6091_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ga0iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6092_o,_al_u6091_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6093|_al_u734  (
    .b({_al_u6002_o,open_n57341}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 }),
    .d({_al_u6092_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [14]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(D*C*~B*~A)"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b0001000000000000),
    .MODE("LOGIC"))
    \_al_u6094|_al_u6889  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ,open_n57362}),
    .b({_al_u6087_o,_al_u6010_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ,_al_u6888_o}),
    .f({_al_u6094_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011000000111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011000000111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6095|_al_u6083  (
    .b({open_n57385,_al_u6082_o}),
    .c({_al_u5998_o,_al_u5998_o}),
    .d({_al_u6079_o,_al_u6079_o}),
    .f({_al_u6095_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6098|_al_u5997  (
    .b({open_n57412,_al_u604_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~B*~(A*~(~D*C)))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0001000100110001),
    .MODE("LOGIC"))
    \_al_u6099|_al_u6097  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ,open_n57433}),
    .b({_al_u6096_o,open_n57434}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 ,_al_u6045_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv }),
    .f({_al_u6099_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6102|_al_u6101  (
    .a({open_n57455,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 }),
    .b({_al_u6101_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6102_o,_al_u6101_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6103|_al_u782  (
    .b({_al_u6002_o,open_n57482}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 }),
    .d({_al_u6102_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6103_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [21]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6106|_al_u6105  (
    .a({open_n57503,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 }),
    .b({_al_u6105_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6106_o,_al_u6105_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6109|_al_u6108  (
    .a({open_n57524,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 }),
    .b({_al_u6108_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6109_o,_al_u6108_o}));
  // ../RTL/cortexm0ds_logic.v(19747)
  EG_PHY_LSLICE #(
    //.LUTF0("~((B*~A)*~(C)*~(D)+(B*~A)*C*~(D)+~((B*~A))*C*D+(B*~A)*C*D)"),
    //.LUTF1("(D*~C*~(~B*~A))"),
    //.LUTG0("~((B*~A)*~(C)*~(D)+(B*~A)*C*~(D)+~((B*~A))*C*D+(B*~A)*C*D)"),
    //.LUTG1("(D*~C*~(~B*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111110111011),
    .INIT_LUTF1(16'b0000111000000000),
    .INIT_LUTG0(16'b0000111110111011),
    .INIT_LUTG1(16'b0000111000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u610|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bi0iu6 ,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0niu6 ,_al_u6989_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u1581_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u609_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jzmiu6 ,open_n57561}),
    .q({open_n57565,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F26bx6 }));  // ../RTL/cortexm0ds_logic.v(19747)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6110|_al_u812  (
    .b({_al_u6006_o,open_n57568}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 }),
    .d({_al_u6109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u6111|_al_u6107  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ,_al_u6002_o}),
    .c({_al_u5998_o,_al_u823_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 ,_al_u6106_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6113|_al_u6112  (
    .a({open_n57615,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 }),
    .b({_al_u6112_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6113_o,_al_u6112_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6114|_al_u794  (
    .b({_al_u6002_o,open_n57642}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 }),
    .d({_al_u6113_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [23]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6116|_al_u6115  (
    .a({open_n57667,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 }),
    .b({_al_u6115_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6116_o,_al_u6115_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*C*B*~A)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*C*B*~A)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6118|_al_u6117  (
    .a({_al_u6104_o,open_n57692}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ,_al_u6002_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ,_al_u6116_o}),
    .f({_al_u6118_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6119|_al_u6916  (
    .b({_al_u6086_o,_al_u6103_o}),
    .c({_al_u6103_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q34ju6_lutinv ,_al_u6915_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M14ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6121|_al_u6120  (
    .a({open_n57739,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 }),
    .b({_al_u6120_o,_al_u823_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6121_o,_al_u6120_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6124|_al_u6123  (
    .a({open_n57760,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 }),
    .b({_al_u6123_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 }),
    .c({_al_u823_o,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6124_o,_al_u6123_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6126|_al_u6125  (
    .a({_al_u6122_o,open_n57781}),
    .b({_al_u6125_o,_al_u6002_o}),
    .c({_al_u6034_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 ,_al_u6124_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T14ju6 ,_al_u6125_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b1000100010100000),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b1000100010100000),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6128|_al_u6127  (
    .a({open_n57806,_al_u6118_o}),
    .b({_al_u6100_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M14ju6 }),
    .c({_al_u6127_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T14ju6 }),
    .d({_al_u6047_o,_al_u5998_o}),
    .f({_al_u6128_o,_al_u6127_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(~A*~(~D*C*~B))"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b0101010101000101),
    .MODE("LOGIC"))
    \_al_u6132|_al_u6130  (
    .a({_al_u6130_o,open_n57831}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ,_al_u604_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u6045_o,_al_u6129_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gy3ju6 ,_al_u6130_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6134|_al_u6133  (
    .a({open_n57852,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 }),
    .b({_al_u6133_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6134_o,_al_u6133_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0101100011111100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0101100011111100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6136|_al_u6026  (
    .a({open_n57877,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .b({_al_u6135_o,_al_u6025_o}),
    .c({_al_u5998_o,_al_u5998_o}),
    .d({_al_u6025_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ,_al_u6026_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6138|_al_u6137  (
    .a({open_n57902,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 }),
    .b({_al_u6137_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6138_o,_al_u6137_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6139|_al_u884  (
    .b({_al_u6002_o,open_n57929}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 }),
    .d({_al_u6138_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({_al_u6139_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [8]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6142|_al_u6141  (
    .a({open_n57950,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 }),
    .b({_al_u6141_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ,_al_u5988_o}),
    .d({_al_u6006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6142_o,_al_u6141_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6143|_al_u890  (
    .b({_al_u6002_o,open_n57973}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 }),
    .d({_al_u6142_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [7]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6145|_al_u6144  (
    .a({open_n57994,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 }),
    .b({_al_u6144_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6145_o,_al_u6144_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*C*~B*~A)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*C*~B*~A)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0001000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6147|_al_u6146  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ,open_n58015}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ,_al_u6006_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ,_al_u6145_o}),
    .f({_al_u6147_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6148|_al_u6140  (
    .b({_al_u6082_o,_al_u6139_o}),
    .c({_al_u6139_o,_al_u5998_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ov3ju6_lutinv ,_al_u6075_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Av3ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u614|_al_u615  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fgpiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6150|_al_u6149  (
    .a({open_n58086,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 }),
    .b({_al_u6149_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6150_o,_al_u6149_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u6152|_al_u6135  (
    .a({_al_u6151_o,open_n58111}),
    .b({_al_u6018_o,_al_u6002_o}),
    .c({_al_u6010_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 }),
    .d({_al_u6135_o,_al_u6134_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu3ju6 ,_al_u6135_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~B*~(~D*~(C*A)))"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b0011001100100000),
    .MODE("LOGIC"))
    \_al_u6154|_al_u6153  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 ,_al_u6147_o}),
    .b({_al_u6128_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Av3ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gy3ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu3ju6 }),
    .d({_al_u6153_o,_al_u5998_o}),
    .f({_al_u6154_o,_al_u6153_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6157|_al_u6156  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .d({_al_u6002_o,_al_u5988_o}),
    .f({_al_u6157_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(~B*A*~(~D*C))"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(~B*A*~(~D*C))"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0010001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6159|_al_u6158  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Queow6 ,open_n58180}),
    .b({_al_u6158_o,_al_u5998_o}),
    .c({_al_u6000_o,_al_u6157_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gweow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .f({_al_u6159_o,_al_u6158_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6161|_al_u6160  (
    .a({open_n58205,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 }),
    .b({_al_u6160_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ,_al_u5988_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1qow6 }),
    .f({_al_u6161_o,_al_u6160_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u6162|_al_u716  (
    .b({_al_u6006_o,open_n58228}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 }),
    .d({_al_u6161_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b0001000100000101),
    .MODE("LOGIC"))
    \_al_u6163|_al_u6151  (
    .a({_al_u6159_o,open_n58249}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 ,_al_u6006_o}),
    .c({_al_u6151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 }),
    .d({_al_u5998_o,_al_u6150_o}),
    .f({_al_u6163_o,_al_u6151_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~A*~(~C*~B)))"),
    //.LUTF1("(B*(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG0("(D*~(~A*~(~C*~B)))"),
    //.LUTG1("(B*(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT_LUTF0(16'b1010101100000000),
    .INIT_LUTF1(16'b1100000001000100),
    .INIT_LUTG0(16'b1010101100000000),
    .INIT_LUTG1(16'b1100000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6166|_al_u6165  (
    .a({_al_u6164_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ,_al_u5998_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ,_al_u5990_o}),
    .d({_al_u6002_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u6166_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0001000100000101),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0001000100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6167|_al_u6025  (
    .a({_al_u6166_o,open_n58294}),
    .b({_al_u6122_o,_al_u6002_o}),
    .c({_al_u6007_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 }),
    .d({_al_u5998_o,_al_u6024_o}),
    .f({_al_u6167_o,_al_u6025_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6168|_al_u6172  (
    .a({open_n58319,_al_u6163_o}),
    .b({open_n58320,_al_u6167_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ,_al_u6169_o}),
    .d({_al_u6164_o,_al_u6171_o}),
    .f({_al_u6168_o,_al_u6172_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(B*~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0100010011000000),
    .MODE("LOGIC"))
    \_al_u6170|_al_u6164  (
    .a({_al_u6164_o,open_n58341}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jbjow6 ,_al_u5998_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv ,_al_u5990_o}),
    .d({_al_u6157_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V2kow6_lutinv }),
    .f({_al_u6170_o,_al_u6164_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*~A)"),
    //.LUTF1("(B*~(~D*~(C*A)))"),
    //.LUTG0("(D*~C*B*~A)"),
    //.LUTG1("(B*~(~D*~(C*A)))"),
    .INIT_LUTF0(16'b0000010000000000),
    .INIT_LUTF1(16'b1100110010000000),
    .INIT_LUTG0(16'b0000010000000000),
    .INIT_LUTG1(16'b1100110010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6173|_al_u6155  (
    .a({_al_u6037_o,_al_u6099_o}),
    .b({_al_u6155_o,_al_u6154_o}),
    .c({_al_u6172_o,_al_u6021_o}),
    .d({_al_u6045_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 }),
    .f({_al_u6173_o,_al_u6155_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u6176|_al_u6175  (
    .a({open_n58386,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u6175_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16]}),
    .d({_al_u2150_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_15 }),
    .f({_al_u6176_o,_al_u6175_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6178|_al_u6174  (
    .a({open_n58407,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 }),
    .b({open_n58408,_al_u1421_o}),
    .c({_al_u6177_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u6174_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 ,_al_u6174_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6181|_al_u6180  (
    .a({open_n58429,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u6180_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ka8ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_10 }),
    .f({_al_u6181_o,_al_u6180_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100000101010),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100000101010),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6183|_al_u6179  (
    .a({open_n58454,_al_u1624_o}),
    .b({open_n58455,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10]}),
    .c({_al_u6182_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I98ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u6183_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I98ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6186|_al_u6185  (
    .a({open_n58480,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u6185_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12]}),
    .d({_al_u2062_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_11 }),
    .f({_al_u6186_o,_al_u6185_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100000101010),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100000101010),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6188|_al_u6184  (
    .a({open_n58505,_al_u1632_o}),
    .b({open_n58506,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 }),
    .c({_al_u6187_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u6184_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u6188_o,_al_u6184_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B*~(C*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000000010011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u6191|_al_u6190  (
    .a({open_n58531,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u6190_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15]}),
    .d({_al_u2128_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_14 }),
    .f({_al_u6191_o,_al_u6190_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100000101010),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6193|_al_u6189  (
    .a({open_n58552,_al_u1413_o}),
    .b({open_n58553,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 }),
    .c({_al_u6192_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u6189_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({_al_u6193_o,_al_u6189_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u6194|_al_u7005  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 ,open_n58574}),
    .b({_al_u6183_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qodow6 }),
    .c({_al_u6188_o,_al_u6980_o}),
    .d({_al_u6193_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 }),
    .f({_al_u6194_o,_al_u7005_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~(D*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0000000100000011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u6197|_al_u6196  (
    .a({open_n58595,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u6196_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[5]}),
    .d({_al_u2252_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24]}),
    .f({_al_u6197_o,_al_u6196_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6199|_al_u6195  (
    .a({open_n58616,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23]}),
    .b({open_n58617,_al_u1485_o}),
    .c({_al_u6198_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Of5ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Of5ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6202|_al_u6201  (
    .a({open_n58638,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u6201_o,_al_u5848_o}),
    .c({_al_u5854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18]}),
    .d({_al_u2171_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_17 }),
    .f({_al_u6202_o,_al_u6201_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100001001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100001001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6204|_al_u6200  (
    .a({open_n58663,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 }),
    .b({open_n58664,_al_u1437_o}),
    .c({_al_u6203_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u6200_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 ,_al_u6200_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~C*~B*~(D*A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000100000011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000100000011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6207|_al_u6206  (
    .a({open_n58689,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 }),
    .b({_al_u6206_o,_al_u5848_o}),
    .c({_al_u5854_o,n1[4]}),
    .d({_al_u2244_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23]}),
    .f({_al_u6207_o,_al_u6206_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000100001001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000100001001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6209|_al_u6205  (
    .a({open_n58714,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 }),
    .b({open_n58715,_al_u1477_o}),
    .c({_al_u6208_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv }),
    .d({_al_u6205_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg5ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 ,_al_u6205_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*D))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000001100001111),
    .INIT_LUT1(16'b1110110101001101),
    .MODE("LOGIC"))
    \_al_u6212|_al_u6211  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [4],open_n58740}),
    .b({_al_u6211_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt4ju6 }),
    .c({_al_u1573_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ys4ju6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wc5ju6_lutinv ,_al_u1573_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl4ju6_lutinv ,_al_u6211_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~B*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6214|_al_u6213  (
    .a({open_n58761,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pk4ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/By4ju6 ,_al_u5848_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_4 }),
    .f({_al_u6214_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4ju6 }));
  // ../RTL/cortexm0ds_logic.v(17907)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~B*~(D*C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0001001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6216|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymzpw6_reg  (
    .a({_al_u5987_o,open_n58786}),
    .b({_al_u6173_o,open_n58787}),
    .c({_al_u6210_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kkkiu6 ,_al_u7041_o}),
    .f({_al_u6216_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .q({open_n58804,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[2] }));  // ../RTL/cortexm0ds_logic.v(17907)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*D))"),
    //.LUTF1("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG0("(~C*~(B*D))"),
    //.LUTG1("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    .INIT_LUTF0(16'b0000001100001111),
    .INIT_LUTF1(16'b1100000011110011),
    .INIT_LUTG0(16'b0000001100001111),
    .INIT_LUTG1(16'b1100000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6217|_al_u2806  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u6216_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv }),
    .f({_al_u6217_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6219|_al_u7095  (
    .c({_al_u6039_o,_al_u6859_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfmow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv }),
    .f({_al_u6219_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*A)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(D*~C*~B*A)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6222|_al_u6220  (
    .a({_al_u6220_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3ju6 ,_al_u6130_o}),
    .c({_al_u6130_o,_al_u6219_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ,_al_u6021_o}),
    .f({_al_u6222_o,_al_u6220_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(~D*A))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0011111100010101),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6223|_al_u6221  (
    .a({open_n58879,_al_u6047_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ,_al_u6050_o}),
    .c({_al_u6219_o,_al_u6087_o}),
    .d({_al_u6222_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3ju6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u6224|_al_u6045  (
    .b({_al_u6044_o,open_n58902}),
    .c({_al_u6041_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 ,_al_u6044_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ,_al_u6045_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b1111101011011101),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b1111101011011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6226|_al_u6104  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ,open_n58923}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ,_al_u6103_o}),
    .c({_al_u6104_o,_al_u5998_o}),
    .d({_al_u6039_o,_al_u6061_o}),
    .f({_al_u6226_o,_al_u6104_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~B*~(~C*A))"),
    //.LUTF1("(C*A*~(~D*B))"),
    //.LUTG0("(D*~B*~(~C*A))"),
    //.LUTG1("(C*A*~(~D*B))"),
    .INIT_LUTF0(16'b0011000100000000),
    .INIT_LUTF1(16'b1010000000100000),
    .INIT_LUTG0(16'b0011000100000000),
    .INIT_LUTG1(16'b1010000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6227|_al_u6225  (
    .a({_al_u6225_o,_al_u6040_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rupow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 }),
    .c({_al_u6226_o,_al_u6035_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u6227_o,_al_u6225_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(~D*~B*~(C*~A))"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000000000100011),
    .MODE("LOGIC"))
    \_al_u6229|_al_u6239  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 ,open_n58972}),
    .b({_al_u6227_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 }),
    .d({_al_u6228_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ru2ju6 }),
    .f({_al_u6229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(~D*~(C*~B))"),
    .INIT_LUT0(16'b0111011100001100),
    .INIT_LUT1(16'b0000000011001111),
    .MODE("LOGIC"))
    \_al_u6231|_al_u6230  (
    .a({open_n58993,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qb3ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M93ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv }),
    .d({_al_u6230_o,_al_u6039_o}),
    .f({_al_u6231_o,_al_u6230_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(B*~(~A*~(D*C)))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b1100100010001000),
    .MODE("LOGIC"))
    \_al_u6233|_al_u6232  (
    .a({_al_u6231_o,open_n59014}),
    .b({_al_u6232_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R83ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u6087_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P73ju6 }),
    .f({_al_u6233_o,_al_u6232_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~((~B*~A))*~(C)+D*(~B*~A)*~(C)+~(D)*(~B*~A)*C+D*(~B*~A)*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("~(D*~((~B*~A))*~(C)+D*(~B*~A)*~(C)+~(D)*(~B*~A)*C+D*(~B*~A)*C)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1110000011101111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1110000011101111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6234|_al_u6236  (
    .a({open_n59035,_al_u6234_o}),
    .b({open_n59036,_al_u6235_o}),
    .c({_al_u6233_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 }),
    .d({_al_u6229_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [33]}),
    .f({_al_u6234_o,_al_u6236_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u6235|_al_u6228  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ,_al_u6044_o}),
    .d({_al_u6228_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7pow6 }),
    .f({_al_u6235_o,_al_u6228_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B@D))"),
    //.LUTF1("(C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    //.LUTG0("(~C*(B@D))"),
    //.LUTG1("(C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    .INIT_LUTF0(16'b0000001100001100),
    .INIT_LUTF1(16'b0010000011100000),
    .INIT_LUTG0(16'b0000001100001100),
    .INIT_LUTG1(16'b0010000011100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6238|_al_u6237  (
    .a({_al_u6236_o,open_n59085}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ng8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .c({_al_u6237_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u6238_o,_al_u6237_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0000001000001110),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b0000001000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6241|_al_u6240  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv ,open_n59110}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fhoiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .c({_al_u6240_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({_al_u6241_o,_al_u6240_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~(D)*~(B)*~(C)+D*~(B)*~(C)+~(D)*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~(D)*~(B)*~(C)+D*~(B)*~(C)+~(D)*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111001111001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6242|_al_u1566  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 ,open_n59137}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32],_al_u1348_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [31],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/To2ju6_lutinv }),
    .f({_al_u6242_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [31]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~B*A*~(D*C))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~B*A*~(D*C))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000001000100010),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6245|_al_u6244  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im2ju6 ,open_n59162}),
    .b({_al_u6244_o,_al_u932_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldoiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u1660_o,_al_u6243_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 ,_al_u6244_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*B*~(C)+D*~(B)*C+~(D)*B*C+D*B*C)"),
    //.LUT1("(C*~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B))"),
    .INIT_LUT0(16'b1111110011000000),
    .INIT_LUT1(16'b0010000011100000),
    .MODE("LOGIC"))
    \_al_u6247|_al_u6246  (
    .a({_al_u6242_o,open_n59187}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .c({_al_u6246_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj2ju6 ,_al_u6246_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~(A)*~(C)*~(D)+A*C*~(D)+A*C*D))"),
    //.LUT1("(~B*~A*~(D@C))"),
    .INIT_LUT0(16'b0010000000100001),
    .INIT_LUT1(16'b0001000000000001),
    .MODE("LOGIC"))
    \_al_u6248|_al_u6218  (
    .a({_al_u6218_o,_al_u6217_o}),
    .b({_al_u6238_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .c({_al_u6241_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj2ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u6248_o,_al_u6218_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6251|_al_u6250  (
    .a({open_n59228,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwiiu6 }),
    .b({_al_u2771_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ai2ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .f({_al_u6251_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ai2ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b1110010011111100),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b1110010011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6254|_al_u6249  (
    .a({_al_u6248_o,open_n59249}),
    .b({_al_u6249_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .c({_al_u6252_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({_al_u6253_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 }),
    .f({_al_u6254_o,_al_u6249_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~B*~A*~(~D*C))"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0001000100000001),
    .MODE("LOGIC"))
    \_al_u6256|_al_u6255  (
    .a({_al_u3208_o,open_n59274}),
    .b({_al_u6255_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N98iu6_lutinv }),
    .c({_al_u1782_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 }),
    .f({_al_u6256_o,_al_u6255_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(C*~B)))"),
    //.LUT1("(A*~(D*C*~B))"),
    .INIT_LUT0(16'b1011101000000000),
    .INIT_LUT1(16'b1000101010101010),
    .MODE("LOGIC"))
    \_al_u6257|_al_u4313  (
    .a({_al_u6256_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv }),
    .b({_al_u1643_o,_al_u1643_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U98iu6 }),
    .d({_al_u1907_o,_al_u1817_o}),
    .f({_al_u6257_o,_al_u4313_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*~(B)*C*D)"),
    //.LUTF1("(A*~(D*~C*~B))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*~(B)*C*D)"),
    //.LUTG1("(A*~(D*~C*~B))"),
    .INIT_LUTF0(16'b0010001111100011),
    .INIT_LUTF1(16'b1010100010101010),
    .INIT_LUTG0(16'b0010001111100011),
    .INIT_LUTG1(16'b1010100010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6260|_al_u6259  (
    .a({_al_u3191_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nsaiu6_lutinv }),
    .b({_al_u6259_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({_al_u606_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .f({_al_u6260_o,_al_u6259_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*~C*B))"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .INIT_LUT0(16'b1010101010100010),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"))
    \_al_u6261|_al_u6258  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yo1ju6 ,_al_u3233_o}),
    .b({_al_u6258_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 }),
    .c({_al_u6260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u6261_o,_al_u6258_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(~D*A))"),
    //.LUTF1("(B*A*~(D*~C))"),
    //.LUTG0("(~(C*B)*~(~D*A))"),
    //.LUTG1("(B*A*~(D*~C))"),
    .INIT_LUTF0(16'b0011111100010101),
    .INIT_LUTF1(16'b1000000010001000),
    .INIT_LUTG0(16'b0011111100010101),
    .INIT_LUTG1(16'b1000000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6263|_al_u6262  (
    .a({_al_u6257_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I82ju6 }),
    .b({_al_u6261_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls1ju6 }),
    .c({_al_u6262_o,_al_u609_o}),
    .d({_al_u3109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u6263_o,_al_u6262_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0101010100000111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0101010100000111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6265|_al_u6266  (
    .a({open_n59383,_al_u3109_o}),
    .b({open_n59384,_al_u6265_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,_al_u2829_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc2ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .f({_al_u6265_o,_al_u6266_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*A))"),
    //.LUTF1("(~D*~C*~(~B*~A))"),
    //.LUTG0("(B*~(D*~C*A))"),
    //.LUTG1("(~D*~C*~(~B*~A))"),
    .INIT_LUTF0(16'b1100010011001100),
    .INIT_LUTF1(16'b0000000000001110),
    .INIT_LUTG0(16'b1100010011001100),
    .INIT_LUTG1(16'b0000000000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6268|_al_u6264  (
    .a({_al_u6264_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eoyiu6_lutinv }),
    .b({_al_u6266_o,_al_u682_o}),
    .c({_al_u6267_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u1907_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u6268_o,_al_u6264_o}));
  // ../RTL/cortexm0ds_logic.v(17512)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(B*A*~(D*~C))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(B*A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110100000101),
    .INIT_LUTF1(16'b1000000010001000),
    .INIT_LUTG0(16'b1111110100000101),
    .INIT_LUTG1(16'b1000000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6269|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6_reg  (
    .a({_al_u6254_o,_al_u6269_o}),
    .b({_al_u6263_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv1ju6 }),
    .c({_al_u6268_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qe8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6269_o,open_n59450}),
    .q({open_n59454,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }));  // ../RTL/cortexm0ds_logic.v(17512)
  // ../RTL/cortexm0ds_logic.v(17765)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b0000000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6271|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7vpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt4iu6 ,open_n59455}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu4iu6 ,open_n59456}),
    .c({_al_u933_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u6271_o,open_n59470}),
    .q({open_n59474,\u_cmsdk_mcu/u_cmsdk_mcu_system/DBGRESTARTED }));  // ../RTL/cortexm0ds_logic.v(17765)
  // ../RTL/cortexm0ds_logic.v(17265)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*A)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(~D*~C*B*A)"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111111111110111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6272|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6_reg  (
    .a({open_n59475,_al_u5643_o}),
    .b({open_n59476,_al_u4452_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u1779_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kt4iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6271_o,_al_u1257_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kt4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt4iu6 }),
    .q({open_n59496,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Isjpw6 }));  // ../RTL/cortexm0ds_logic.v(17265)
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(D*~A*~(~C*~B))"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(D*~A*~(~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0101010000000000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0101010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6280|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b3  (
    .a({_al_u6276_o,\u_cmsdk_mcu/HADDR [10]}),
    .b({_al_u6277_o,\u_cmsdk_mcu/HADDR [4]}),
    .c({_al_u6278_o,\u_cmsdk_mcu/HADDR [3]}),
    .clk(XTAL1_wire),
    .d({_al_u6279_o,\u_cmsdk_mcu/HADDR [2]}),
    .mi({open_n59501,\u_cmsdk_mcu/HADDR [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6280_o,_al_u6278_o}),
    .q({open_n59516,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(D*C*~B*A)"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"))
    \_al_u6289|_al_u6290  (
    .a({_al_u4921_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 ,_al_u6289_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }),
    .f({_al_u6289_o,_al_u6290_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u6292|_al_u6291  (
    .a({_al_u4551_o,_al_u4091_o}),
    .b({_al_u6291_o,_al_u4101_o}),
    .c({_al_u4035_o,_al_u4126_o}),
    .d({_al_u4086_o,_al_u4131_o}),
    .f({_al_u6292_o,_al_u6291_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*~A)"),
    //.LUT1("(B*A*~(~D*~C))"),
    .INIT_LUT0(16'b0100000000000000),
    .INIT_LUT1(16'b1000100010000000),
    .MODE("LOGIC"))
    \_al_u6294|_al_u6293  (
    .a({\u_cmsdk_mcu/HADDR [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xg6iu6 }),
    .b({\u_cmsdk_mcu/HSIZE [1],_al_u4919_o}),
    .c({_al_u6290_o,_al_u6292_o}),
    .d({_al_u6293_o,_al_u4056_o}),
    .f({_al_u6294_o,_al_u6293_o}));
  // ../RTL/cortexm0ds_logic.v(17670)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~A*~(~C*~B))"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110101011),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6304|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6_reg  (
    .a({open_n59577,_al_u6295_o}),
    .b({open_n59578,_al_u5000_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 ,\u_cmsdk_mcu/HADDR [8]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u6304_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6304_o,open_n59592}),
    .q({open_n59596,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzspw6 }));  // ../RTL/cortexm0ds_logic.v(17670)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6307|_al_u6308  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wh0ju6 ,open_n59597}),
    .b({_al_u4376_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 ,_al_u6307_o}),
    .f({_al_u6307_o,_al_u6308_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*~C*~A))"),
    //.LUT1("(~C*~(B*~D))"),
    .INIT_LUT0(16'b1100110011001000),
    .INIT_LUT1(16'b0000111100000011),
    .MODE("LOGIC"))
    \_al_u6310|_al_u6309  (
    .a({open_n59622,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6ziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwjax6 }),
    .d({_al_u6308_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .f({_al_u6310_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T6ziu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~B*(C@A))"),
    //.LUTF1("(C*~(~B*~D))"),
    //.LUTG0("(~D*~B*(C@A))"),
    //.LUTG1("(C*~(~B*~D))"),
    .INIT_LUTF0(16'b0000000000010010),
    .INIT_LUTF1(16'b1111000011000000),
    .INIT_LUTG0(16'b0000000000010010),
    .INIT_LUTG1(16'b1111000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6311|_al_u6306  (
    .a({open_n59643,_al_u6248_o}),
    .b({_al_u6310_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6ziu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0piu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({_al_u6306_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 }),
    .f({_al_u6311_o,_al_u6306_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~D*~B*~(C*~A))"),
    //.LUTG0("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*~(C)*D+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~D*~B*~(C*~A))"),
    .INIT_LUTF0(16'b1010100000101000),
    .INIT_LUTF1(16'b0000000000100011),
    .INIT_LUTG0(16'b1010100000101000),
    .INIT_LUTG1(16'b0000000000100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6314|_al_u6313  (
    .a({_al_u6313_o,_al_u6312_o}),
    .b({_al_u3419_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4kax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P14qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4jax6 }),
    .f({_al_u6314_o,_al_u6313_o}));
  // ../RTL/cortexm0ds_logic.v(17240)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*~A))"),
    //.LUTF1("(D*~(~A*~(~C*B)))"),
    //.LUTG0("(~(~D*C)*~(B*~A))"),
    //.LUTG1("(D*~(~A*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b1010111000000000),
    .INIT_LUTG0(16'b1011101100001011),
    .INIT_LUTG1(16'b1010111000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6315|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6_reg  (
    .a({_al_u6311_o,_al_u6315_o}),
    .b({_al_u3183_o,_al_u6329_o}),
    .c({_al_u6314_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u2868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }),
    .f({_al_u6315_o,open_n59710}),
    .q({open_n59714,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgjpw6 }));  // ../RTL/cortexm0ds_logic.v(17240)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~D*C*~B*~A)"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~D*C*~B*~A)"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000010000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6317|_al_u6316  (
    .a({_al_u1784_o,_al_u3223_o}),
    .b({_al_u1801_o,_al_u1367_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeziu6 ,_al_u3124_o}),
    .d({_al_u6316_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .f({_al_u6317_o,_al_u6316_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~A*~(D*C*B))"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"))
    \_al_u6321|_al_u6320  (
    .a({_al_u6320_o,_al_u903_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv ,_al_u3094_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6kiu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u1266_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvjpw6 }),
    .f({_al_u6321_o,_al_u6320_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6322|_al_u6319  (
    .b({_al_u6319_o,_al_u4161_o}),
    .c({_al_u6321_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u3664_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z37ow6_lutinv }),
    .f({_al_u6322_o,_al_u6319_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6323|_al_u4414  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxyiu6 ,open_n59787}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gebow6_lutinv ,_al_u1775_o}),
    .d({_al_u6322_o,_al_u3109_o}),
    .f({_al_u6323_o,_al_u4414_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~C*~(~D*B*A))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000111100000111),
    .MODE("LOGIC"))
    \_al_u6325|_al_u6324  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuyiu6_lutinv ,open_n59808}),
    .b({_al_u4393_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .c({_al_u6324_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sojax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ssjax6 ,_al_u2364_o}),
    .f({_al_u6325_o,_al_u6324_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(~D*C))"),
    //.LUT1("(B*A*~(~D*C))"),
    .INIT_LUT0(16'b1000100000001000),
    .INIT_LUT1(16'b1000100000001000),
    .MODE("LOGIC"))
    \_al_u6326|_al_u6318  (
    .a({_al_u6318_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Veziu6 }),
    .b({_al_u6323_o,_al_u6317_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htyiu6 ,_al_u3202_o}),
    .d({_al_u6325_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dxvpw6 }),
    .f({_al_u6326_o,_al_u6318_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*~A*~(D*B))"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000100000101),
    .MODE("LOGIC"))
    \_al_u6327|_al_u3568  (
    .a({_al_u3101_o,open_n59849}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3ziu6 ,_al_u1271_o}),
    .c({_al_u3236_o,_al_u1342_o}),
    .d({_al_u1271_o,_al_u1266_o}),
    .f({_al_u6327_o,_al_u3568_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(~D*~C))"),
    //.LUTF1("(~C*A*~(D*B))"),
    //.LUTG0("(B*A*~(~D*~C))"),
    //.LUTG1("(~C*A*~(D*B))"),
    .INIT_LUTF0(16'b1000100010000000),
    .INIT_LUTF1(16'b0000001000001010),
    .INIT_LUTG0(16'b1000100010000000),
    .INIT_LUTG1(16'b0000001000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6328|_al_u6329  (
    .a({_al_u6327_o,_al_u6326_o}),
    .b({_al_u2361_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcziu6 }),
    .c({_al_u3078_o,_al_u6328_o}),
    .d({_al_u3401_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 }),
    .f({_al_u6328_o,_al_u6329_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*~A*~(~D*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*~A*~(~D*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0101000000010000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0101000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6331|_al_u5330  (
    .a({_al_u5329_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ,_al_u927_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ,_al_u5329_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 }),
    .f({_al_u6331_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogqiu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(C*~(~B*D))"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6333|_al_u6332  (
    .a({open_n59918,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 }),
    .b({_al_u6332_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 }),
    .d({_al_u6331_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 }),
    .f({_al_u6333_o,_al_u6332_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6335|_al_u3375  (
    .a({open_n59943,_al_u2725_o}),
    .b({open_n59944,_al_u1301_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ch5iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 }),
    .f({_al_u6335_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ag5iu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6337|_al_u6338  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nt9bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C10bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 }),
    .f({_al_u6337_o,_al_u6338_o}));
  // ../RTL/cortexm0ds_logic.v(20087)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*B*~(~C*A))"),
    //.LUT1("(B*~(~C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6340|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6_reg  (
    .a({open_n59997,_al_u6337_o}),
    .b({_al_u6338_o,_al_u6338_o}),
    .c({_al_u6339_o,_al_u6339_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6337_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 }),
    .mi({open_n60008,\u_cmsdk_mcu/HWDATA [22]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 ,_al_u6350_o}),
    .q({open_n60012,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 }));  // ../RTL/cortexm0ds_logic.v(20087)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6342|_al_u573  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [1]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Czzax6 ,_al_u470_o}),
    .f({_al_u6342_o,_al_u573_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6343|_al_u6354  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ikhbx6 ,_al_u6343_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 ,_al_u6342_o}),
    .f({_al_u6343_o,_al_u6354_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(B*~(~C*A)))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0000000000111011),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u6345|_al_u6347  (
    .a({open_n60065,_al_u6342_o}),
    .b({_al_u6343_o,_al_u6343_o}),
    .c({_al_u6344_o,_al_u6344_o}),
    .d({_al_u6342_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 }),
    .f({_al_u6345_o,_al_u6347_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6346|_al_u5300  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 }),
    .d({_al_u6345_o,_al_u5299_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv ,_al_u5300_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(B)*~((~C*A))*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+~(B)*(~C*A)*D)"),
    //.LUTF1("(~D*B*~(~C*A))"),
    //.LUTG0("(~(B)*~((~C*A))*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+~(B)*(~C*A)*D)"),
    //.LUTG1("(~D*B*~(~C*A))"),
    .INIT_LUTF0(16'b1111011100110001),
    .INIT_LUTF1(16'b0000000011000100),
    .INIT_LUTG0(16'b1111011100110001),
    .INIT_LUTG1(16'b0000000011000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6348|_al_u6344  (
    .a({_al_u6342_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 }),
    .b({_al_u6343_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 }),
    .c({_al_u6344_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yryax6 }),
    .f({_al_u6348_o,_al_u6344_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    //.LUT1("(~D*~(B*~(~C*A)))"),
    .INIT_LUT0(16'b1101010011110101),
    .INIT_LUT1(16'b0000000000111011),
    .MODE("LOGIC"))
    \_al_u6349|_al_u6339  (
    .a({_al_u6337_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 }),
    .b({_al_u6338_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 }),
    .c({_al_u6339_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cwyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tngbx6 }),
    .f({_al_u6349_o,_al_u6339_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6352|_al_u6341  (
    .b({open_n60158,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 }),
    .c({_al_u6338_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eyyax6 }),
    .d({_al_u6337_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 }),
    .f({_al_u6352_o,_al_u6341_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~((~D*~A))+~B*C*~((~D*~A))+~(~B)*C*(~D*~A)+~B*C*(~D*~A))"),
    //.LUTF1("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    //.LUTG0("(~B*~(C)*~((~D*~A))+~B*C*~((~D*~A))+~(~B)*C*(~D*~A)+~B*C*(~D*~A))"),
    //.LUTG1("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT_LUTF0(16'b0011001101110010),
    .INIT_LUTF1(16'b0000000011101000),
    .INIT_LUTG0(16'b0011001101110010),
    .INIT_LUTG1(16'b0000000011101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6353|_al_u6355  (
    .a({_al_u6341_o,_al_u6353_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv ,_al_u6341_o}),
    .c({_al_u6351_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oltow6_lutinv }),
    .d({_al_u6352_o,_al_u6354_o}),
    .f({_al_u6353_o,_al_u6355_o}));
  // ../RTL/cortexm0ds_logic.v(19107)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6356|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ,open_n60203}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 }),
    .mi({open_n60207,\u_cmsdk_mcu/HWDATA [31]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6356_o,_al_u6361_o}),
    .q({open_n60222,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 }));  // ../RTL/cortexm0ds_logic.v(19107)
  // ../RTL/cortexm0ds_logic.v(19113)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(C*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6359|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6_reg  (
    .b({_al_u6357_o,_al_u6358_o}),
    .c({_al_u6358_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6356_o,_al_u6357_o}),
    .mi({open_n60228,\u_cmsdk_mcu/HWDATA [30]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ,_al_u6369_o}),
    .q({open_n60243,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uizax6 }));  // ../RTL/cortexm0ds_logic.v(19113)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(~D*C))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1000100000001000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6360|_al_u6357  (
    .a({open_n60244,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owhbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgzax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 }),
    .f({_al_u6360_o,_al_u6357_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6362|_al_u5659  (
    .b({open_n60267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U31bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C3wpw6 ,_al_u5658_o}),
    .f({_al_u6362_o,_al_u5659_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6365|_al_u6366  (
    .b({_al_u6363_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 }),
    .c({_al_u6364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 }),
    .d({_al_u6362_o,_al_u6365_o}),
    .f({_al_u6365_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~D*A*~(C*~B))"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~D*A*~(C*~B))"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b0000000010001010),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b0000000010001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6368|_al_u6363  (
    .a({_al_u6362_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 }),
    .b({_al_u6363_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 }),
    .c({_al_u6364_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 }),
    .f({_al_u6368_o,_al_u6363_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~D*C*~(B*~A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000010110000),
    .MODE("LOGIC"))
    \_al_u6370|_al_u5153  (
    .a({_al_u6356_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 }),
    .b({_al_u6357_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 }),
    .c({_al_u6358_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 }),
    .f({_al_u6370_o,_al_u5153_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~B*D))"),
    //.LUTF1("(~B*~A*~(~D*~C))"),
    //.LUTG0("(~C*~(~B*D))"),
    //.LUTG1("(~B*~A*~(~D*~C))"),
    .INIT_LUTF0(16'b0000110000001111),
    .INIT_LUTF1(16'b0001000100010000),
    .INIT_LUTG0(16'b0000110000001111),
    .INIT_LUTG1(16'b0001000100010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6371|_al_u6367  (
    .a({_al_u6367_o,open_n60358}),
    .b({_al_u6368_o,_al_u6364_o}),
    .c({_al_u6369_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 }),
    .d({_al_u6370_o,_al_u6362_o}),
    .f({_al_u6371_o,_al_u6367_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~((~D*~A))+~B*C*~((~D*~A))+~(~B)*C*(~D*~A)+~B*C*(~D*~A))"),
    //.LUTF1("(~A*(B*C*~(D)+B*~(C)*D+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~B*~(C)*~((~D*~A))+~B*C*~((~D*~A))+~(~B)*C*(~D*~A)+~B*C*(~D*~A))"),
    //.LUTG1("(~A*(B*C*~(D)+B*~(C)*D+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0011001101110010),
    .INIT_LUTF1(16'b0101010001000000),
    .INIT_LUTG0(16'b0011001101110010),
    .INIT_LUTG1(16'b0101010001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6372|_al_u6374  (
    .a({_al_u6360_o,_al_u6372_o}),
    .b({_al_u6361_o,_al_u6361_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttow6_lutinv }),
    .d({_al_u6371_o,_al_u6373_o}),
    .f({_al_u6372_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(~D*C))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1000100000001000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6373|_al_u6364  (
    .a({open_n60407,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aa2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cxzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 }),
    .d({_al_u6362_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 }),
    .f({_al_u6373_o,_al_u6364_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111000011100100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6375|_al_u6377  (
    .a({open_n60428,_al_u6353_o}),
    .b({open_n60429,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjtow6_lutinv }),
    .c({_al_u6348_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjtow6_lutinv }),
    .d({_al_u6347_o,_al_u6354_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjtow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(~D*~C))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~B*~A*~(~D*~C))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0001000100010000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0001000100010000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6376|_al_u6351  (
    .a({open_n60450,_al_u6347_o}),
    .b({open_n60451,_al_u6348_o}),
    .c({_al_u6350_o,_al_u6349_o}),
    .d({_al_u6349_o,_al_u6350_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjtow6_lutinv ,_al_u6351_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6378|_al_u6384  (
    .c({_al_u6368_o,_al_u6373_o}),
    .d({_al_u6367_o,_al_u6360_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwtow6_lutinv ,_al_u6384_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6379|_al_u6358  (
    .c({_al_u6370_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5bbx6 }),
    .d({_al_u6369_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1bbx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tktow6_lutinv ,_al_u6358_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*A)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(D*~C*~B*A)"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u637|_al_u596  (
    .a({open_n60528,_al_u379_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full }),
    .f({_al_u637_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n61 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111000011100100),
    .MODE("LOGIC"))
    \_al_u6380|_al_u6601  (
    .a({_al_u6372_o,open_n60553}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iwtow6_lutinv ,_al_u6372_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tktow6_lutinv ,_al_u6373_o}),
    .d({_al_u6373_o,_al_u6385_o}),
    .f({_al_u6380_o,_al_u6601_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*~(B*~A)))"),
    //.LUT1("(~(D*~C)*~(B*~A))"),
    .INIT_LUT0(16'b1111000001000000),
    .INIT_LUT1(16'b1011000010111011),
    .MODE("LOGIC"))
    \_al_u6381|_al_u6437  (
    .a({_al_u6355_o,_al_u6381_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ,_al_u6383_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8tow6_lutinv }),
    .d({_al_u6380_o,_al_u6384_o}),
    .f({_al_u6381_o,_al_u6437_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6382|_al_u6647  (
    .c({_al_u6354_o,_al_u6354_o}),
    .d({_al_u6352_o,_al_u6353_o}),
    .f({_al_u6382_o,_al_u6647_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~C*~(~B*D))"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000110000001111),
    .MODE("LOGIC"))
    \_al_u6383|_al_u6386  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv ,_al_u6355_o}),
    .c({_al_u6382_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oetow6_lutinv }),
    .d({_al_u6355_o,_al_u6385_o}),
    .f({_al_u6383_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~(B*~A))"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(~D*C*~(B*~A))"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b0000000010110000),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000000010110000),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6385|_al_u6438  (
    .a({open_n60640,_al_u6381_o}),
    .b({_al_u6383_o,_al_u6383_o}),
    .c({_al_u6384_o,_al_u6380_o}),
    .d({_al_u6381_o,_al_u6384_o}),
    .f({_al_u6385_o,_al_u6438_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6387|_al_u6388  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fc1bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D70bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C50bx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ,_al_u6388_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(A)*~((C*~B))*~(D)+~(A)*~((C*~B))*D+A*~((C*~B))*D+~(A)*(C*~B)*D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1101111101000101),
    .MODE("LOGIC"))
    \_al_u6389|_al_u5029  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 }),
    .f({_al_u6389_o,_al_u5029_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6392|_al_u6393  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkjbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Us3bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rijbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C30bx6 }),
    .f({_al_u6392_o,_al_u6393_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*B*~(~C*A))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(~D*B*~(~C*A))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011000100),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000000011000100),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6395|_al_u6398  (
    .a({open_n60737,_al_u6392_o}),
    .b({_al_u6393_o,_al_u6393_o}),
    .c({_al_u6394_o,_al_u6394_o}),
    .d({_al_u6392_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 }),
    .f({_al_u6395_o,_al_u6398_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    //.LUTF1("(~D*~(B*~(~C*A)))"),
    //.LUTG0("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    //.LUTG1("(~D*~(B*~(~C*A)))"),
    .INIT_LUTF0(16'b1101010011110101),
    .INIT_LUTF1(16'b0000000000111011),
    .INIT_LUTG0(16'b1101010011110101),
    .INIT_LUTG1(16'b0000000000111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6397|_al_u6394  (
    .a({_al_u6392_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 }),
    .b({_al_u6393_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 }),
    .c({_al_u6394_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 }),
    .f({_al_u6397_o,_al_u6394_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6402|_al_u6390  (
    .b({open_n60788,_al_u6388_o}),
    .c({_al_u6388_o,_al_u6389_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 }),
    .f({_al_u6402_o,_al_u6390_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~((~D*~A))+B*C*~((~D*~A))+~(B)*C*(~D*~A)+B*C*(~D*~A))"),
    //.LUTF1("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    //.LUTG0("(B*~(C)*~((~D*~A))+B*C*~((~D*~A))+~(B)*C*(~D*~A)+B*C*(~D*~A))"),
    //.LUTG1("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    .INIT_LUTF0(16'b1100110011011000),
    .INIT_LUTF1(16'b0000000010110010),
    .INIT_LUTG0(16'b1100110011011000),
    .INIT_LUTG1(16'b0000000010110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6403|_al_u6405  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv ,_al_u6403_o}),
    .b({_al_u6396_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv }),
    .c({_al_u6401_o,_al_u6396_o}),
    .d({_al_u6402_o,_al_u6404_o}),
    .f({_al_u6403_o,_al_u6405_o}));
  // ../RTL/cortexm0ds_logic.v(19197)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6406|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6_reg  (
    .a({open_n60833,\u_cmsdk_mcu/HWDATA [13]}),
    .b({open_n60834,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6406_o,open_n60848}),
    .q({open_n60852,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 }));  // ../RTL/cortexm0ds_logic.v(19197)
  // ../RTL/cortexm0ds_logic.v(19191)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000011111000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0111000011111000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6407|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6_reg  (
    .a({open_n60853,\u_cmsdk_mcu/HWDATA [12]}),
    .b({open_n60854,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6407_o,open_n60872}),
    .q({open_n60876,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90bx6 }));  // ../RTL/cortexm0ds_logic.v(19191)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1101010011110101),
    .MODE("LOGIC"))
    \_al_u6408|_al_u6713  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 }),
    .f({_al_u6408_o,_al_u6713_o}));
  // ../RTL/cortexm0ds_logic.v(19873)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*B*~(~C*A))"),
    //.LUT1("(B*~(~C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6409|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6_reg  (
    .a({open_n60897,_al_u6406_o}),
    .b({_al_u6407_o,_al_u6407_o}),
    .c({_al_u6408_o,_al_u6408_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6406_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 }),
    .mi({open_n60908,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6409_o,_al_u6417_o}),
    .q({open_n60912,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7abx6 }));  // ../RTL/cortexm0ds_logic.v(19873)
  // ../RTL/cortexm0ds_logic.v(19209)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110001000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1101111110001000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6411|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6_reg  (
    .a({open_n60913,\u_cmsdk_mcu/HWDATA [15]}),
    .b({open_n60914,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V59iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6411_o,open_n60932}),
    .q({open_n60936,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 }));  // ../RTL/cortexm0ds_logic.v(19209)
  // ../RTL/cortexm0ds_logic.v(19203)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6412|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6_reg  (
    .a({open_n60937,\u_cmsdk_mcu/HWDATA [14]}),
    .b({open_n60938,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6412_o,open_n60952}),
    .q({open_n60956,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 }));  // ../RTL/cortexm0ds_logic.v(19203)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1101010011110101),
    .MODE("LOGIC"))
    \_al_u6413|_al_u5154  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 }),
    .f({_al_u6413_o,_al_u5154_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*B*~(~C*A))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0000000011000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u6414|_al_u6419  (
    .a({open_n60977,_al_u6411_o}),
    .b({_al_u6412_o,_al_u6412_o}),
    .c({_al_u6413_o,_al_u6413_o}),
    .d({_al_u6411_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pjgbx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 ,_al_u6419_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(B*~(~C*A)))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000000111011),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6421|_al_u6418  (
    .a({open_n60998,_al_u6411_o}),
    .b({open_n60999,_al_u6412_o}),
    .c({_al_u6412_o,_al_u6413_o}),
    .d({_al_u6411_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M85bx6 }),
    .f({_al_u6421_o,_al_u6418_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    //.LUT1("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b1111000010110001),
    .INIT_LUT1(16'b0000000011101000),
    .MODE("LOGIC"))
    \_al_u6422|_al_u6424  (
    .a({_al_u6410_o,_al_u6422_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv ,_al_u6410_o}),
    .c({_al_u6420_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv }),
    .d({_al_u6421_o,_al_u6423_o}),
    .f({_al_u6422_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B*~(~C*A)))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~(B*~(~C*A)))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000111011),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000111011),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6423|_al_u6416  (
    .a({open_n61040,_al_u6406_o}),
    .b({open_n61041,_al_u6407_o}),
    .c({_al_u6407_o,_al_u6408_o}),
    .d({_al_u6406_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G25bx6 }),
    .f({_al_u6423_o,_al_u6416_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000011100100),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000011100100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6425|_al_u6427  (
    .a({open_n61066,_al_u6403_o}),
    .b({open_n61067,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Akuow6_lutinv }),
    .c({_al_u6398_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8uow6_lutinv }),
    .d({_al_u6397_o,_al_u6404_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Akuow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(~D*~C))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0001000100010000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6426|_al_u6401  (
    .a({open_n61092,_al_u6397_o}),
    .b({open_n61093,_al_u6398_o}),
    .c({_al_u6400_o,_al_u6399_o}),
    .d({_al_u6399_o,_al_u6400_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8uow6_lutinv ,_al_u6401_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~((~D*~A))+C*B*~((~D*~A))+~(C)*B*(~D*~A)+C*B*(~D*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111000011100100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6428|_al_u6430  (
    .a({open_n61114,_al_u6422_o}),
    .b({open_n61115,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7uow6_lutinv }),
    .c({_al_u6417_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8uow6_lutinv }),
    .d({_al_u6416_o,_al_u6423_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7uow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(~D*~C))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0001000100010000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6429|_al_u6420  (
    .a({open_n61136,_al_u6416_o}),
    .b({open_n61137,_al_u6417_o}),
    .c({_al_u6419_o,_al_u6418_o}),
    .d({_al_u6418_o,_al_u6419_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8uow6_lutinv ,_al_u6420_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(~D*C)*~(B*~A))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(~D*C)*~(B*~A))"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1011101100001011),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1011101100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6431|_al_u6436  (
    .a({_al_u6405_o,open_n61158}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv ,_al_u6405_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv ,_al_u6435_o}),
    .f({_al_u6431_o,_al_u6436_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6434|_al_u6404  (
    .c({_al_u6402_o,_al_u6393_o}),
    .d({_al_u6404_o,_al_u6392_o}),
    .f({_al_u6434_o,_al_u6404_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~B*D))"),
    //.LUT1("(~B*~(~C*~D))"),
    .INIT_LUT0(16'b0000110000001111),
    .INIT_LUT1(16'b0011001100110000),
    .MODE("LOGIC"))
    \_al_u6439|_al_u6433  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3uow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdtow6_lutinv }),
    .c({_al_u6434_o,_al_u6432_o}),
    .d({_al_u6433_o,_al_u6405_o}),
    .f({_al_u6439_o,_al_u6433_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(~D*~C*~(B*~A))"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(~D*~C*~(B*~A))"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b0000000000001011),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0000000000001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6440|_al_u6435  (
    .a({_al_u6431_o,open_n61229}),
    .b({_al_u6433_o,_al_u6433_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yctow6_lutinv ,_al_u6434_o}),
    .d({_al_u6434_o,_al_u6431_o}),
    .f({_al_u6440_o,_al_u6435_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6442|_al_u6446  (
    .b({open_n61256,_al_u6435_o}),
    .c({_al_u6432_o,_al_u6432_o}),
    .d({_al_u6435_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 }),
    .f({_al_u6442_o,_al_u6446_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    //.LUT1("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b0000111101001110),
    .INIT_LUT1(16'b0000000011101000),
    .MODE("LOGIC"))
    \_al_u6443|_al_u6556  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv ,_al_u6443_o}),
    .b({_al_u6436_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irrow6_lutinv }),
    .c({_al_u6441_o,_al_u6436_o}),
    .d({_al_u6442_o,_al_u6444_o}),
    .f({_al_u6443_o,_al_u6556_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6444|_al_u6445  (
    .c({_al_u6382_o,_al_u6444_o}),
    .d({_al_u6384_o,_al_u6443_o}),
    .f({_al_u6444_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6447|_al_u5305  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9abx6 }),
    .f({_al_u6447_o,_al_u5305_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTF1("(B*A*~(D*~C))"),
    //.LUTG0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG1("(B*A*~(D*~C))"),
    .INIT_LUTF0(16'b0000110011111100),
    .INIT_LUTF1(16'b1000000010001000),
    .INIT_LUTG0(16'b0000110011111100),
    .INIT_LUTG1(16'b1000000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6448|_al_u2743  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 ,open_n61349}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 ,\u_cmsdk_mcu/sram_hrdata [29]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ,\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ,_al_u2741_o}),
    .f({_al_u6448_o,\u_cmsdk_mcu/u_ahb_ram/n13 [29]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~(B*~A))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b0000000010110000),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u6450|_al_u6458  (
    .a({open_n61374,_al_u6447_o}),
    .b({_al_u6448_o,_al_u6448_o}),
    .c({_al_u6449_o,_al_u6449_o}),
    .d({_al_u6447_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 }),
    .f({_al_u6450_o,_al_u6458_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"))
    \_al_u6451|_al_u6464  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bc3bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kojpw6 }),
    .d({_al_u6450_o,_al_u6450_o}),
    .f({_al_u6451_o,_al_u6464_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6455|_al_u6459  (
    .b({_al_u6453_o,_al_u6454_o}),
    .c({_al_u6454_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 }),
    .d({_al_u6452_o,_al_u6453_o}),
    .f({_al_u6455_o,_al_u6459_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~D*C*~(B*~A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~D*C*~(B*~A))"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b0000000010110000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b0000000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6460|_al_u6452  (
    .a({_al_u6452_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 }),
    .b({_al_u6453_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 }),
    .c({_al_u6454_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 }),
    .f({_al_u6460_o,_al_u6452_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(~B*~A*~(~D*~C))"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(~B*~A*~(~D*~C))"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b0001000100010000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0001000100010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6461|_al_u6457  (
    .a({_al_u6457_o,open_n61467}),
    .b({_al_u6458_o,_al_u6449_o}),
    .c({_al_u6459_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Up4bx6 }),
    .d({_al_u6460_o,_al_u6448_o}),
    .f({_al_u6461_o,_al_u6457_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~(~D*A))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(C*B*~(~D*A))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1100000001000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000001000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6462|_al_u6453  (
    .a({open_n61492,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hg3bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S0kbx6 }),
    .d({_al_u6455_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 ,_al_u6453_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(B)*~((~C*~A))+~D*B*~((~C*~A))+~(~D)*B*(~C*~A)+~D*B*(~C*~A))"),
    //.LUT1("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b1111101100000001),
    .INIT_LUT1(16'b0000000011101000),
    .MODE("LOGIC"))
    \_al_u6463|_al_u6465  (
    .a({_al_u6451_o,_al_u6463_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv ,_al_u6451_o}),
    .c({_al_u6461_o,_al_u6464_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmrow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv }),
    .f({_al_u6463_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6467|_al_u3502  (
    .b({open_n61539,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5upw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jz2bx6 ,_al_u2725_o}),
    .f({_al_u6467_o,_al_u3502_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(A)*~(C)*~((D*~B))+~(A)*C*~((D*~B))+A*C*~((D*~B))+~(A)*C*(D*~B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1101010011110101),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1101010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6468|_al_u6806  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 }),
    .f({_al_u6468_o,_al_u6806_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*B*~(~C*A))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(~D*B*~(~C*A))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011000100),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000000011000100),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6469|_al_u6479  (
    .a({open_n61588,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 }),
    .b({_al_u6467_o,_al_u6467_o}),
    .c({_al_u6468_o,_al_u6468_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 }),
    .f({_al_u6469_o,_al_u6479_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6473|_al_u3491  (
    .b({open_n61615,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oxkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv2bx6 ,_al_u2717_o}),
    .f({_al_u6473_o,_al_u3491_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~D))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b0000111100000011),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u6474|_al_u6476  (
    .b({_al_u6472_o,_al_u6473_o}),
    .c({_al_u6473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 }),
    .d({_al_u6471_o,_al_u6472_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ,_al_u6476_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~D*C*~(B*~A))"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b0000000010110000),
    .MODE("LOGIC"))
    \_al_u6477|_al_u6471  (
    .a({_al_u6471_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 }),
    .b({_al_u6472_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 }),
    .c({_al_u6473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 }),
    .f({_al_u6477_o,_al_u6471_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~A*~(~D*~C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~A*~(~D*~C))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001000100010000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001000100010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6480|_al_u6466  (
    .a({_al_u6476_o,open_n61678}),
    .b({_al_u6477_o,open_n61679}),
    .c({_al_u6478_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qx0bx6 }),
    .d({_al_u6479_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P33bx6 }),
    .f({_al_u6480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B*~(~C*A)))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~(B*~(~C*A)))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000111011),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000111011),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6481|_al_u6478  (
    .a({open_n61704,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 }),
    .b({open_n61705,_al_u6467_o}),
    .c({_al_u6467_o,_al_u6468_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amsow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E34bx6 }),
    .f({_al_u6481_o,_al_u6478_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000010110010),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000010110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6482|_al_u6475  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv ,open_n61730}),
    .b({_al_u6475_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 }),
    .c({_al_u6480_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 }),
    .d({_al_u6481_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 }),
    .f({_al_u6482_o,_al_u6475_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~(~D*A))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(C*B*~(~D*A))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1100000001000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100000001000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6483|_al_u6472  (
    .a({open_n61755,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv0bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rm2bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wu3bx6 }),
    .f({_al_u6483_o,_al_u6472_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1111000111100000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1111000111100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6484|_al_u6613  (
    .a({_al_u6482_o,open_n61780}),
    .b({_al_u6483_o,_al_u6482_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv ,_al_u6483_o}),
    .d({_al_u6475_o,_al_u6495_o}),
    .f({_al_u6484_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111111000010000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111111000010000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6485|_al_u6487  (
    .a({open_n61805,_al_u6482_o}),
    .b({open_n61806,_al_u6483_o}),
    .c({_al_u6477_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqsow6_lutinv }),
    .d({_al_u6476_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqsow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqsow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6486|_al_u6494  (
    .c({_al_u6479_o,_al_u6481_o}),
    .d({_al_u6478_o,_al_u6483_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pqsow6_lutinv ,_al_u6494_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111111000010000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111111000010000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6488|_al_u6490  (
    .a({open_n61859,_al_u6463_o}),
    .b({open_n61860,_al_u6464_o}),
    .c({_al_u6458_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzsow6_lutinv }),
    .d({_al_u6457_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzsow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzsow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6489|_al_u6454  (
    .c({_al_u6460_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcipw6 }),
    .d({_al_u6459_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz0bx6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzsow6_lutinv ,_al_u6454_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(~D*C)*~(~B*A))"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1101110100001101),
    .MODE("LOGIC"))
    \_al_u6491|_al_u6496  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv ,open_n61909}),
    .b({_al_u6484_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv ,_al_u6484_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv ,_al_u6495_o}),
    .f({_al_u6491_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6497|_al_u5040  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 }),
    .f({_al_u6497_o,_al_u5040_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6499|_al_u5203  (
    .b({open_n61956,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P12bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hbpow6_lutinv }),
    .f({_al_u6499_o,_al_u5203_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~(B*~A))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b0000000010110000),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u6500|_al_u6508  (
    .a({open_n61981,_al_u6497_o}),
    .b({_al_u6498_o,_al_u6498_o}),
    .c({_al_u6499_o,_al_u6499_o}),
    .d({_al_u6497_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhgbx6 }),
    .f({_al_u6500_o,_al_u6508_o}));
  // ../RTL/cortexm0ds_logic.v(19221)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTF1("(C*A*~(D*~B))"),
    //.LUTG0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTG1("(C*A*~(D*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000011111000),
    .INIT_LUTF1(16'b1000000010100000),
    .INIT_LUTG0(16'b0111000011111000),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6503|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ,\u_cmsdk_mcu/HWDATA [17]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6503_o,open_n62019}),
    .q({open_n62023,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 }));  // ../RTL/cortexm0ds_logic.v(19221)
  // ../RTL/cortexm0ds_logic.v(19215)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111000011111000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6504|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6_reg  (
    .a({open_n62024,\u_cmsdk_mcu/HWDATA [16]}),
    .b({open_n62025,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6504_o,open_n62039}),
    .q({open_n62043,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 }));  // ../RTL/cortexm0ds_logic.v(19215)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~D))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b0000111100000011),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u6505|_al_u6509  (
    .b({_al_u6503_o,_al_u6504_o}),
    .c({_al_u6504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 }),
    .d({_al_u6502_o,_al_u6503_o}),
    .f({_al_u6505_o,_al_u6509_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6506|_al_u6515  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 }),
    .d({_al_u6505_o,_al_u6505_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv ,_al_u6515_o}));
  // ../RTL/cmsdk_apb_uart.v(592)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*~D))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("~(~B*~(C*~D))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011111100),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1100110011111100),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u650|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ,open_n62092}),
    .b({_al_u473_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample }),
    .c({_al_u467_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n106 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0],_al_u650_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u650_o,open_n62109}),
    .q({open_n62113,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full }));  // ../RTL/cmsdk_apb_uart.v(592)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~D*C*~(B*~A))"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b0000000010110000),
    .MODE("LOGIC"))
    \_al_u6510|_al_u6502  (
    .a({_al_u6502_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 }),
    .b({_al_u6503_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 }),
    .c({_al_u6504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5abx6 }),
    .f({_al_u6510_o,_al_u6502_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(~D*~C*~(~B*~A))"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(~D*~C*~(~B*~A))"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b0000000000001110),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0000000000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6511|_al_u6507  (
    .a({_al_u6507_o,open_n62134}),
    .b({_al_u6508_o,_al_u6499_o}),
    .c({_al_u6509_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pczax6 }),
    .d({_al_u6510_o,_al_u6498_o}),
    .f({_al_u6511_o,_al_u6507_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*A*~(C*~B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1000101000000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6512|_al_u6498  (
    .a({open_n62159,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ln0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 }),
    .d({_al_u6500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V52bx6 }),
    .f({_al_u6512_o,_al_u6498_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    //.LUTF1("(~D*(~(A)*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C))"),
    //.LUTG0("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    //.LUTG1("(~D*(~(A)*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT_LUTF0(16'b1111000111100000),
    .INIT_LUTF1(16'b0000000011010100),
    .INIT_LUTG0(16'b1111000111100000),
    .INIT_LUTG1(16'b0000000011010100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6513|_al_u6539  (
    .a({_al_u6501_o,_al_u6513_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv ,_al_u6515_o}),
    .c({_al_u6511_o,_al_u6501_o}),
    .d({_al_u6512_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J2sow6_lutinv }),
    .f({_al_u6513_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~((~C*~A))+B*D*~((~C*~A))+~(B)*D*(~C*~A)+B*D*(~C*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100110111001000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6514|_al_u6517  (
    .a({open_n62204,_al_u6513_o}),
    .b({open_n62205,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3sow6_lutinv }),
    .c({_al_u6508_o,_al_u6515_o}),
    .d({_al_u6507_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L3sow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3sow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(19251)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTF1("(D*A*~(C*~B))"),
    //.LUTG0("~(~C*~(D)*~((B*A))+~C*D*~((B*A))+~(~C)*D*(B*A)+~C*D*(B*A))"),
    //.LUTG1("(D*A*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000011111000),
    .INIT_LUTF1(16'b1000101000000000),
    .INIT_LUTG0(16'b0111000011111000),
    .INIT_LUTG1(16'b1000101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6519|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ,\u_cmsdk_mcu/HWDATA [23]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O59iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6519_o,open_n62243}),
    .q({open_n62247,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 }));  // ../RTL/cortexm0ds_logic.v(19251)
  // ../RTL/cortexm0ds_logic.v(19023)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~D))"),
    //.LUT1("(C*~(B*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000011),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6521|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6_reg  (
    .b({_al_u6519_o,_al_u6520_o}),
    .c({_al_u6520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6518_o,_al_u6519_o}),
    .mi({open_n62260,\u_cmsdk_mcu/HWDATA [30]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6521_o,_al_u6529_o}),
    .q({open_n62264,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 }));  // ../RTL/cortexm0ds_logic.v(19023)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6522|_al_u6803  (
    .a({open_n62265,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ot0bx6 }),
    .d({_al_u6521_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xq2bx6 }),
    .f({_al_u6522_o,_al_u6803_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(C*A*~(D*~B))"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b1000000010100000),
    .MODE("LOGIC"))
    \_al_u6525|_al_u3476  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 ,open_n62286}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ,\u_cmsdk_mcu/HWDATA [21]}),
    .f({_al_u6525_o,_al_u3476_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6527|_al_u6531  (
    .b({_al_u6525_o,_al_u6526_o}),
    .c({_al_u6526_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 }),
    .d({_al_u6524_o,_al_u6525_o}),
    .f({_al_u6527_o,_al_u6531_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~D*C*~(B*~A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~D*C*~(B*~A))"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b0000000010110000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b0000000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6530|_al_u6518  (
    .a({_al_u6518_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 }),
    .b({_al_u6519_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 }),
    .c({_al_u6520_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Unyax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 }),
    .f({_al_u6530_o,_al_u6518_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~D*C*~(B*~A))"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~D*C*~(B*~A))"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b0000000010110000),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b0000000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6532|_al_u6524  (
    .a({_al_u6524_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 }),
    .b({_al_u6525_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 }),
    .c({_al_u6526_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 }),
    .f({_al_u6532_o,_al_u6524_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    //.LUTF1("(~A*(~(B)*C*~(D)+~(B)*~(C)*D+~(B)*C*D+B*C*D))"),
    //.LUTG0("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    //.LUTG1("(~A*(~(B)*C*~(D)+~(B)*~(C)*D+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b1111000111100000),
    .INIT_LUTF1(16'b0101000100010000),
    .INIT_LUTG0(16'b1111000111100000),
    .INIT_LUTG1(16'b0101000100010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6534|_al_u6540  (
    .a({_al_u6522_o,_al_u6534_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv ,_al_u6535_o}),
    .c({_al_u6528_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv }),
    .d({_al_u6533_o,_al_u6528_o}),
    .f({_al_u6534_o,_al_u6540_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*~(D)*~((~B*~A))+C*D*~((~B*~A))+~(C)*D*(~B*~A)+C*D*(~B*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000111100000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000111100000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6536|_al_u6538  (
    .a({open_n62405,_al_u6534_o}),
    .b({open_n62406,_al_u6535_o}),
    .c({_al_u6530_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6sow6_lutinv }),
    .d({_al_u6529_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3sow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D6sow6_lutinv ,_al_u6538_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~(~B*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~C*~(~B*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001110),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001110),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6537|_al_u6533  (
    .a({open_n62431,_al_u6529_o}),
    .b({open_n62432,_al_u6530_o}),
    .c({_al_u6532_o,_al_u6531_o}),
    .d({_al_u6531_o,_al_u6532_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3sow6_lutinv ,_al_u6533_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~(B*~A))"),
    //.LUTF1("(~(~D*C)*~(~B*A))"),
    //.LUTG0("(~D*C*~(B*~A))"),
    //.LUTG1("(~(~D*C)*~(~B*A))"),
    .INIT_LUTF0(16'b0000000010110000),
    .INIT_LUTF1(16'b1101110100001101),
    .INIT_LUTG0(16'b0000000010110000),
    .INIT_LUTG1(16'b1101110100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6541|_al_u6547  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv ,_al_u6541_o}),
    .b({_al_u6538_o,_al_u6543_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ewrow6_lutinv }),
    .d({_al_u6540_o,_al_u6544_o}),
    .f({_al_u6541_o,_al_u6547_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6542|_al_u6523  (
    .b({open_n62483,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 }),
    .c({_al_u6535_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpyax6 }),
    .d({_al_u6522_o,_al_u6521_o}),
    .f({_al_u6542_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1sow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6544|_al_u6620  (
    .c({_al_u6512_o,_al_u6515_o}),
    .d({_al_u6515_o,_al_u6513_o}),
    .f({_al_u6544_o,_al_u6620_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*~(B*~A)))"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(C*~(~D*~(B*~A)))"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b1111000001000000),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b1111000001000000),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6545|_al_u6548  (
    .a({open_n62528,_al_u6541_o}),
    .b({_al_u6543_o,_al_u6543_o}),
    .c({_al_u6544_o,_al_u6538_o}),
    .d({_al_u6541_o,_al_u6544_o}),
    .f({_al_u6545_o,_al_u6548_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6546|_al_u6639  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv ,open_n62555}),
    .c({_al_u6540_o,_al_u6545_o}),
    .d({_al_u6545_o,_al_u6558_o}),
    .f({_al_u6546_o,_al_u6639_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~C)*~(~B*~A))"),
    //.LUTF1("(~B*~(~C*~D))"),
    //.LUTG0("(~(~D*~C)*~(~B*~A))"),
    //.LUTG1("(~B*~(~C*~D))"),
    .INIT_LUTF0(16'b1110111011100000),
    .INIT_LUTF1(16'b0011001100110000),
    .INIT_LUTG0(16'b1110111011100000),
    .INIT_LUTG1(16'b0011001100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6549|_al_u6551  (
    .a({open_n62580,_al_u6547_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rksow6_lutinv ,_al_u6548_o}),
    .c({_al_u6494_o,_al_u6549_o}),
    .d({_al_u6493_o,_al_u6550_o}),
    .f({_al_u6549_o,_al_u6551_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~D))"),
    //.LUT1("(~D*~C*~(B*~A))"),
    .INIT_LUT0(16'b0000111100000011),
    .INIT_LUT1(16'b0000000000001011),
    .MODE("LOGIC"))
    \_al_u6550|_al_u6495  (
    .a({_al_u6491_o,open_n62605}),
    .b({_al_u6493_o,_al_u6493_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yksow6_lutinv ,_al_u6494_o}),
    .d({_al_u6494_o,_al_u6491_o}),
    .f({_al_u6550_o,_al_u6495_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~D))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000111100000011),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6552|_al_u6493  (
    .b({open_n62628,_al_u6484_o}),
    .c({_al_u6492_o,_al_u6492_o}),
    .d({_al_u6495_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxrow6_lutinv }),
    .f({_al_u6552_o,_al_u6493_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(~D*(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b0000000011101000),
    .MODE("LOGIC"))
    \_al_u6553|_al_u6570  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv ,open_n62649}),
    .b({_al_u6546_o,_al_u6558_o}),
    .c({_al_u6551_o,_al_u6552_o}),
    .d({_al_u6552_o,_al_u6446_o}),
    .f({_al_u6553_o,_al_u6570_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~D))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000111100000011),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6554|_al_u6543  (
    .b({open_n62672,_al_u6540_o}),
    .c({_al_u6542_o,_al_u6542_o}),
    .d({_al_u6545_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxrow6_lutinv }),
    .f({_al_u6554_o,_al_u6543_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(~B*~(D)*~((~C*~A))+~B*D*~((~C*~A))+~(~B)*D*(~C*~A)+~B*D*(~C*~A))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100100011001101),
    .MODE("LOGIC"))
    \_al_u6555|_al_u6558  (
    .a({_al_u6553_o,open_n62693}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gqrow6_lutinv ,open_n62694}),
    .c({_al_u6554_o,_al_u6554_o}),
    .d({_al_u6546_o,_al_u6553_o}),
    .f({_al_u6555_o,_al_u6558_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6557|_al_u6567  (
    .b({open_n62717,_al_u6555_o}),
    .c({_al_u6556_o,_al_u6556_o}),
    .d({_al_u6555_o,_al_u6566_o}),
    .f({_al_u6557_o,_al_u6567_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000101000011111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000101000011111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6559|_al_u6560  (
    .a({open_n62742,_al_u6553_o}),
    .b({open_n62743,_al_u6554_o}),
    .c({_al_u6550_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mtrow6_lutinv }),
    .d({_al_u6549_o,_al_u6547_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mtrow6_lutinv ,_al_u6560_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000111101001110),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6561|_al_u6563  (
    .a({open_n62768,_al_u6443_o}),
    .b({open_n62769,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kctow6_lutinv }),
    .c({_al_u6438_o,_al_u6562_o}),
    .d({_al_u6437_o,_al_u6444_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kctow6_lutinv ,_al_u6563_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~C)*~(~B*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(~D*~C)*~(~B*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1110111011100000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1110111011100000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6562|_al_u6441  (
    .a({open_n62790,_al_u6437_o}),
    .b({open_n62791,_al_u6438_o}),
    .c({_al_u6440_o,_al_u6439_o}),
    .d({_al_u6439_o,_al_u6440_o}),
    .f({_al_u6562_o,_al_u6441_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(D*~A))"),
    //.LUT1("(~A*~(D*~(~C*~B)))"),
    .INIT_LUT0(16'b1010100011111100),
    .INIT_LUT1(16'b0000000101010101),
    .MODE("LOGIC"))
    \_al_u6566|_al_u6565  (
    .a({_al_u6446_o,_al_u6558_o}),
    .b({_al_u6557_o,_al_u6555_o}),
    .c({_al_u6564_o,_al_u6556_o}),
    .d({_al_u6565_o,_al_u6552_o}),
    .f({_al_u6566_o,_al_u6565_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~(D*A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~C*B*~(D*A))"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0000010000001100),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000010000001100),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6568|_al_u6564  (
    .a({open_n62836,_al_u6558_o}),
    .b({_al_u6560_o,_al_u6560_o}),
    .c({_al_u6548_o,_al_u6563_o}),
    .d({_al_u6558_o,_al_u6548_o}),
    .f({_al_u6568_o,_al_u6564_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~((C*~A))+B*D*~((C*~A))+~(B)*D*(C*~A)+B*D*(C*~A))"),
    //.LUTF1("(~C*(~(A)*B*~(D)+~(A)*~(B)*D+~(A)*B*D+A*B*D))"),
    //.LUTG0("(B*~(D)*~((C*~A))+B*D*~((C*~A))+~(B)*D*(C*~A)+B*D*(C*~A))"),
    //.LUTG1("(~C*(~(A)*B*~(D)+~(A)*~(B)*D+~(A)*B*D+A*B*D))"),
    .INIT_LUTF0(16'b1101110010001100),
    .INIT_LUTF1(16'b0000110100000100),
    .INIT_LUTG0(16'b1101110010001100),
    .INIT_LUTG1(16'b0000110100000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6571|_al_u6574  (
    .a({_al_u6567_o,_al_u6571_o}),
    .b({_al_u6569_o,_al_u6567_o}),
    .c({_al_u6570_o,_al_u6572_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 }),
    .f({_al_u6571_o,_al_u6574_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6572|_al_u5093  (
    .b({open_n62887,_al_u5067_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdtpw6 }),
    .d({_al_u5329_o,_al_u5092_o}),
    .f({_al_u6572_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~((C*~A))+B*D*~((C*~A))+~(B)*D*(C*~A)+B*D*(C*~A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(D)*~((C*~A))+B*D*~((C*~A))+~(B)*D*(C*~A)+B*D*(C*~A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1101110010001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1101110010001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6573|_al_u6580  (
    .a({open_n62908,_al_u6571_o}),
    .b({open_n62909,_al_u6579_o}),
    .c({_al_u6572_o,_al_u6572_o}),
    .d({_al_u6571_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 }),
    .f({_al_u6573_o,_al_u6580_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6575|_al_u927  (
    .c({_al_u5329_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnwiu6 }),
    .d({_al_u6570_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuciu6 }),
    .f({_al_u6575_o,_al_u927_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~D*~(B*~A)))"),
    //.LUT1("(~(~D*B)*~(~C*~A))"),
    .INIT_LUT0(16'b0000111100000100),
    .INIT_LUT1(16'b1111101000110010),
    .MODE("LOGIC"))
    \_al_u6576|_al_u6599  (
    .a({_al_u6573_o,_al_u6582_o}),
    .b({_al_u6574_o,_al_u6576_o}),
    .c({_al_u6575_o,_al_u6573_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ,_al_u6335_o}),
    .f({_al_u6576_o,_al_u6599_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u6578|_al_u6577  (
    .b({_al_u6577_o,open_n62984}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ,_al_u6574_o}),
    .d({_al_u6336_o,_al_u6576_o}),
    .f({_al_u6578_o,_al_u6577_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b1110010000000000),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"))
    \_al_u6579|_al_u6569  (
    .a({open_n63005,_al_u6566_o}),
    .b({_al_u6568_o,_al_u6568_o}),
    .c({_al_u6563_o,_al_u6563_o}),
    .d({_al_u6566_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wgipw6 }),
    .f({_al_u6579_o,_al_u6569_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(~D*~B)*~(C*~A))"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b1010111110001100),
    .MODE("LOGIC"))
    \_al_u6582|_al_u6581  (
    .a({_al_u6574_o,open_n63026}),
    .b({_al_u6580_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 }),
    .d({_al_u6581_o,_al_u6333_o}),
    .f({_al_u6582_o,_al_u6581_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~(B*~A))"),
    //.LUT1("(C*~(~D*~(B*~A)))"),
    .INIT_LUT0(16'b0000000000001011),
    .INIT_LUT1(16'b1111000001000000),
    .MODE("LOGIC"))
    \_al_u6584|_al_u6583  (
    .a({_al_u6582_o,_al_u6582_o}),
    .b({_al_u6576_o,_al_u6576_o}),
    .c({_al_u6580_o,_al_u6333_o}),
    .d({_al_u6335_o,_al_u6335_o}),
    .f({_al_u6584_o,_al_u6583_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~(C*~B)))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .INIT_LUT0(16'b0010000010101010),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"))
    \_al_u6586|_al_u6636  (
    .a({_al_u6582_o,_al_u6631_o}),
    .b({_al_u6576_o,_al_u6582_o}),
    .c({_al_u3722_o,_al_u6576_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ffrow6_lutinv ,_al_u6333_o}),
    .f({_al_u6586_o,_al_u6636_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~A*~(D*~B))"),
    //.LUTF1("(~D*~(~C*~(~B*~A)))"),
    //.LUTG0("(~C*~A*~(D*~B))"),
    //.LUTG1("(~D*~(~C*~(~B*~A)))"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000000011110001),
    .INIT_LUTG0(16'b0000010000000101),
    .INIT_LUTG1(16'b0000000011110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6588|_al_u4264  (
    .a({_al_u6336_o,_al_u4261_o}),
    .b({_al_u6577_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0biu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sbrow6 ,_al_u4263_o}),
    .d({_al_u3749_o,_al_u3753_o}),
    .f({_al_u6588_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li5iu6 }));
  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u658|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b6  (
    .b({open_n63113,_al_u569_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n7_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux9_b10_sel_is_3_o ,open_n63130}),
    .q({open_n63134,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [6]}));  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~D))"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0011001100000011),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u6590|_al_u6589  (
    .b({_al_u6575_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F17ax6 }),
    .c({_al_u6589_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnmpw6 }),
    .d({_al_u6573_o,_al_u5329_o}),
    .f({_al_u6590_o,_al_u6589_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~(~B*A)))"),
    //.LUT1("(D*~(C*~(B*~A)))"),
    .INIT_LUT0(16'b1111001000000000),
    .INIT_LUT1(16'b0100111100000000),
    .MODE("LOGIC"))
    \_al_u6592|_al_u6795  (
    .a({_al_u6578_o,_al_u6592_o}),
    .b({_al_u6587_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv }),
    .c({_al_u6588_o,_al_u6593_o}),
    .d({_al_u6591_o,_al_u5067_o}),
    .f({_al_u6592_o,_al_u6795_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~B*~(~C*~(D*~A)))"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0011000100110000),
    .MODE("LOGIC"))
    \_al_u6593|_al_u1791  (
    .a({_al_u1774_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M8row6_lutinv }),
    .b({_al_u1791_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A9row6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }),
    .f({_al_u6593_o,_al_u1791_o}));
  // ../RTL/cortexm0ds_logic.v(18589)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*C)*~(~B*~A))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100010001),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6595|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xfiax6_reg  (
    .a({open_n63197,_al_u1882_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oy8iu6 ,_al_u1906_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stuow6_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n590 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cz8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iixpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oy8iu6 }),
    .q({open_n63213,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_primask_o }));  // ../RTL/cortexm0ds_logic.v(18589)
  // ../RTL/cortexm0ds_logic.v(17468)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*~(~B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000110000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6596|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6_reg  (
    .a({open_n63214,_al_u6592_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K7row6_lutinv ,_al_u6593_o}),
    .c({_al_u6593_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u6592_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6596_o,open_n63228}),
    .q({open_n63232,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 }));  // ../RTL/cortexm0ds_logic.v(17468)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6597|_al_u1386  (
    .b({_al_u1385_o,open_n63235}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnnpw6 ,_al_u1385_o}),
    .d({_al_u2855_o,_al_u1299_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3row6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/HALTED }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6600|_al_u6611  (
    .c({_al_u6566_o,_al_u6566_o}),
    .d({_al_u6599_o,_al_u6599_o}),
    .f({_al_u6600_o,_al_u6611_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    //.LUT1("~(~B*~((D*~C))*~(A)+~B*(D*~C)*~(A)+~(~B)*(D*~C)*A+~B*(D*~C)*A)"),
    .INIT_LUT0(16'b0000101000011111),
    .INIT_LUT1(16'b1110010011101110),
    .MODE("LOGIC"))
    \_al_u6603|_al_u6602  (
    .a({_al_u6385_o,_al_u6353_o}),
    .b({_al_u6602_o,_al_u6354_o}),
    .c({_al_u6372_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hkgow6 }),
    .d({_al_u6365_o,_al_u6345_o}),
    .f({_al_u6603_o,_al_u6602_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6604|_al_u6609  (
    .b({_al_u6603_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfgow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjgow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gggow6_lutinv }),
    .d({_al_u6601_o,_al_u6435_o}),
    .f({_al_u6604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6605|_al_u6410  (
    .b({open_n63332,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E05bx6 }),
    .c({_al_u6423_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 }),
    .d({_al_u6422_o,_al_u6409_o}),
    .f({_al_u6605_o,_al_u6410_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6606|_al_u6415  (
    .b({_al_u6409_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa5bx6 }),
    .d({_al_u6605_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whgow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfgow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G9uow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6607|_al_u6391  (
    .b({open_n63381,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 }),
    .c({_al_u6404_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sh4bx6 }),
    .d({_al_u6403_o,_al_u6390_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phuow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u6608|_al_u6396  (
    .b({_al_u6390_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 }),
    .c({_al_u6395_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 ,_al_u6395_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gggow6_lutinv ,_al_u6396_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b0010101000001000),
    .MODE("LOGIC"))
    \_al_u6610|_al_u6634  (
    .a({_al_u6600_o,_al_u6600_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 }),
    .c({_al_u6604_o,_al_u6435_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgow6_lutinv ,_al_u6385_o}),
    .f({_al_u6610_o,_al_u6634_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~(D*A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0001000000110000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6612|_al_u6587  (
    .a({open_n63448,_al_u6583_o}),
    .b({open_n63449,_al_u6584_o}),
    .c({_al_u6590_o,_al_u6586_o}),
    .d({_al_u6583_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vpgbx6 }),
    .f({_al_u6612_o,_al_u6587_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6614|_al_u6618  (
    .c({_al_u6464_o,_al_u6614_o}),
    .d({_al_u6463_o,_al_u6495_o}),
    .f({_al_u6614_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6615|_al_u6470  (
    .b({open_n63500,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odgow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G54bx6 }),
    .d({_al_u6482_o,_al_u6469_o}),
    .f({_al_u6615_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Upsow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C)*~(A)+~(~D*B)*C*~(A)+~(~(~D*B))*C*A+~(~D*B)*C*A)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~(~D*B)*~(C)*~(A)+~(~D*B)*C*~(A)+~(~(~D*B))*C*A+~(~D*B)*C*A)"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b1111010110110001),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111010110110001),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6617|_al_u6616  (
    .a({open_n63521,_al_u6495_o}),
    .b({_al_u6616_o,_al_u6614_o}),
    .c({_al_u6469_o,_al_u6615_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv ,_al_u6450_o}),
    .f({_al_u6617_o,_al_u6616_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6619|_al_u6456  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cy4bx6 }),
    .c({_al_u6455_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 }),
    .d({_al_u6617_o,_al_u6455_o}),
    .f({_al_u6619_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpsow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6621|_al_u6501  (
    .b({_al_u6500_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 }),
    .c({_al_u6505_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rezax6 }),
    .d({_al_u6620_o,_al_u6500_o}),
    .f({_al_u6621_o,_al_u6501_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000101000011111),
    .MODE("LOGIC"))
    \_al_u6622|_al_u6535  (
    .a({_al_u6534_o,open_n63598}),
    .b({_al_u6535_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li2bx6 }),
    .c({_al_u6521_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr0bx6 }),
    .d({_al_u6527_o,_al_u6527_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pagow6_lutinv ,_al_u6535_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0000111111001100),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u6625|_al_u6624  (
    .a({_al_u6610_o,open_n63619}),
    .b({_al_u6611_o,_al_u6619_o}),
    .c({_al_u6612_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bagow6_lutinv }),
    .d({_al_u6624_o,_al_u6558_o}),
    .f({_al_u6625_o,_al_u6624_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~B*~(~C*~D))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~B*~(~C*~D))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011001100110000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011001100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6626|_al_u5380  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 ,_al_u5067_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T8kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyax6 }),
    .d({_al_u6625_o,_al_u5379_o}),
    .f({_al_u6626_o,_al_u5380_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u6627|_al_u6775  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ,_al_u6745_o}),
    .d({_al_u6626_o,_al_u6655_o}),
    .f({_al_u6627_o,_al_u6775_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C@B)*~(D@A))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1000001001000001),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6629|_al_u6638  (
    .a({open_n63690,_al_u6633_o}),
    .b({open_n63691,_al_u6637_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 }),
    .d({_al_u6600_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 }),
    .f({_al_u6629_o,_al_u6638_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B*~A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(D*~(~C*~B*~A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1111111000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111111000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6631|_al_u6649  (
    .a({open_n63712,_al_u6643_o}),
    .b({open_n63713,_al_u6648_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv ,_al_u6590_o}),
    .d({_al_u6590_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0fow6_lutinv }),
    .f({_al_u6631_o,_al_u6649_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6632|_al_u5149  (
    .b({_al_u6631_o,_al_u5143_o}),
    .c({_al_u6558_o,_al_u5148_o}),
    .d({_al_u6611_o,_al_u5067_o}),
    .f({_al_u6632_o,_al_u5149_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*B*~A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b1011000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6633|_al_u6695  (
    .a({open_n63764,_al_u6629_o}),
    .b({open_n63765,_al_u6632_o}),
    .c({_al_u6632_o,_al_u6694_o}),
    .d({_al_u6629_o,_al_u5067_o}),
    .f({_al_u6633_o,_al_u6695_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6637|_al_u6635  (
    .a({open_n63786,_al_u6611_o}),
    .b({_al_u6635_o,_al_u6558_o}),
    .c({_al_u6636_o,_al_u6495_o}),
    .d({_al_u6634_o,_al_u6545_o}),
    .f({_al_u6637_o,_al_u6635_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0011001111110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u6640|_al_u6623  (
    .b({open_n63813,_al_u6621_o}),
    .c({_al_u6620_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pagow6_lutinv }),
    .d({_al_u6545_o,_al_u6545_o}),
    .f({_al_u6640_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bagow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    //.LUT1("(~B*~(A*~(~D*~C)))"),
    .INIT_LUT0(16'b1111111001010100),
    .INIT_LUT1(16'b0001000100010011),
    .MODE("LOGIC"))
    \_al_u6642|_al_u6641  (
    .a({_al_u6639_o,_al_u6558_o}),
    .b({_al_u6641_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C8fow6 }),
    .c({_al_u6534_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8fow6_lutinv }),
    .d({_al_u6535_o,_al_u6640_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1fow6 ,_al_u6641_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6643|_al_u6591  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1fow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0biu6 }),
    .d({_al_u6611_o,_al_u6590_o}),
    .f({_al_u6643_o,_al_u6591_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6646|_al_u6645  (
    .b({_al_u6601_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4fow6 }),
    .c({_al_u6645_o,_al_u6605_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 ,_al_u6435_o}),
    .f({_al_u6646_o,_al_u6645_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*A*~(~D*B))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*A*~(~D*B))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000101000000010),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000101000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6648|_al_u6644  (
    .a({_al_u6600_o,open_n63904}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2fow6 ,open_n63905}),
    .c({_al_u6646_o,_al_u6385_o}),
    .d({_al_u6647_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4fow6 }),
    .f({_al_u6648_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2fow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~(D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*B*~(D*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000010000001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000010000001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6650|_al_u3541  (
    .a({open_n63930,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Am7ow6 }),
    .b({open_n63931,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kubow6 }),
    .c({_al_u6631_o,_al_u3540_o}),
    .d({_al_u6600_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 }),
    .f({_al_u6650_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtbow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6652|_al_u6661  (
    .b({open_n63958,_al_u6660_o}),
    .c({_al_u6631_o,_al_u5067_o}),
    .d({_al_u6611_o,_al_u6652_o}),
    .f({_al_u6652_o,_al_u6661_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*D))"),
    //.LUTF1("(~(C@B)*~(D*~A))"),
    //.LUTG0("(C*~(~B*D))"),
    //.LUTG1("(~(C@B)*~(D*~A))"),
    .INIT_LUTF0(16'b1100000011110000),
    .INIT_LUTF1(16'b1000001011000011),
    .INIT_LUTG0(16'b1100000011110000),
    .INIT_LUTG1(16'b1000001011000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6653|_al_u6651  (
    .a({_al_u6650_o,open_n63983}),
    .b({_al_u6652_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ,_al_u6650_o}),
    .f({_al_u6653_o,_al_u6651_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*(D@A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0100000010000000),
    .MODE("LOGIC"))
    \_al_u6654|_al_u3248  (
    .a({_al_u6649_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc8iu6 }),
    .b({_al_u6651_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Habiu6 }),
    .c({_al_u6653_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .f({_al_u6654_o,_al_u3248_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(D*C*~A))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1000110011001100),
    .MODE("LOGIC"))
    \_al_u6655|_al_u6628  (
    .a({_al_u6627_o,open_n64028}),
    .b({_al_u6628_o,open_n64029}),
    .c({_al_u6638_o,_al_u1299_o}),
    .d({_al_u6654_o,_al_u6596_o}),
    .f({_al_u6655_o,_al_u6628_o}));
  // ../RTL/cortexm0ds_logic.v(17284)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(D*C*~B))"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("~(~A*~(D*C*~B))"),
    //.LUTG1("(~C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010101010),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1011101010101010),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6656|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6_reg  (
    .a({open_n64050,_al_u6655_o}),
    .b({_al_u1777_o,_al_u6656_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,_al_u1299_o}),
    .clk(XTAL1_wire),
    .d({_al_u6596_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6656_o,open_n64068}),
    .q({open_n64072,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }));  // ../RTL/cortexm0ds_logic.v(17284)
  // ../RTL/cortexm0ds_logic.v(17709)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6659|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,open_n64073}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,_al_u2173_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 ,_al_u2171_o}),
    .f({_al_u6659_o,\u_cmsdk_mcu/HWDATA [17]}),
    .q({open_n64094,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjupw6 }));  // ../RTL/cortexm0ds_logic.v(17709)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u6660|_al_u6658  (
    .a({_al_u6658_o,open_n64095}),
    .b({_al_u6659_o,_al_u5260_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jj0bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dt1bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }),
    .f({_al_u6660_o,_al_u6658_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*A*~(D*B))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0010000010100000),
    .MODE("LOGIC"))
    \_al_u6664|_al_u6662  (
    .a({_al_u6662_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .c({_al_u6663_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Erbbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 }),
    .f({_al_u6664_o,_al_u6662_o}));
  // ../RTL/cortexm0ds_logic.v(20212)
  EG_PHY_LSLICE #(
    //.LUTF0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTF1("(~D*A*~(C*~B))"),
    //.LUTG0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTG1("(~D*A*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000100000001),
    .INIT_LUTF1(16'b0000000010001010),
    .INIT_LUTG0(16'b1111000100000001),
    .INIT_LUTG1(16'b0000000010001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6668|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6_reg  (
    .a({_al_u6666_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({_al_u1833_o,_al_u1833_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({_al_u6667_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 }),
    .f({_al_u6668_o,open_n64154}),
    .q({open_n64158,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tujbx6 }));  // ../RTL/cortexm0ds_logic.v(20212)
  // ../RTL/cortexm0ds_logic.v(19930)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~B*~(D*A))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111001111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6670|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6_reg  (
    .a({open_n64159,_al_u5053_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u6669_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 ,_al_u6670_o}),
    .clk(XTAL1_wire),
    .d({_al_u5049_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yubbx6 }),
    .f({_al_u6670_o,open_n64174}),
    .q({open_n64178,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 }));  // ../RTL/cortexm0ds_logic.v(19930)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6673|_al_u6672  (
    .a({open_n64179,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .b({_al_u3779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }),
    .c({_al_u5260_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ih0bx6 }),
    .d({_al_u6672_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jx1bx6 }),
    .f({_al_u6673_o,_al_u6672_o}));
  // ../RTL/cortexm0ds_logic.v(17658)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6674|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,open_n64204}),
    .b({_al_u405_o,_al_u2290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T2kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 ,_al_u2289_o}),
    .f({_al_u6674_o,\u_cmsdk_mcu/HWDATA [16]}),
    .q({open_n64225,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujspw6 }));  // ../RTL/cortexm0ds_logic.v(17658)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u6676|_al_u6683  (
    .b({_al_u6675_o,_al_u6676_o}),
    .c({_al_u5067_o,_al_u6682_o}),
    .d({_al_u6650_o,_al_u5020_o}),
    .f({_al_u6676_o,_al_u6683_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u6679|_al_u6678  (
    .a({_al_u6677_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjtiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owcax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 }),
    .f({_al_u6679_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjtiu6 }));
  // ../RTL/cortexm0ds_logic.v(18183)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6680|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,_al_u4049_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4048_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Chwpw6 }),
    .mi({open_n64278,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .f({_al_u6680_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dbmiu6 }),
    .q({open_n64283,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kcaax6 }));  // ../RTL/cortexm0ds_logic.v(18183)
  // ../RTL/cortexm0ds_logic.v(18317)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6681|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6_reg  (
    .a({_al_u6679_o,open_n64284}),
    .b({_al_u6680_o,open_n64285}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .mi({open_n64296,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .f({_al_u6681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 }),
    .q({open_n64301,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aoeax6 }));  // ../RTL/cortexm0ds_logic.v(18317)
  // ../RTL/cortexm0ds_logic.v(18647)
  EG_PHY_MSLICE #(
    //.LUT0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUT1("(~D*A*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100000001),
    .INIT_LUT1(16'b0000000010001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6682|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6_reg  (
    .a({_al_u6681_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({_al_u1868_o,_al_u1868_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .clk(XTAL1_wire),
    .d({_al_u6667_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 }),
    .f({_al_u6682_o,open_n64316}),
    .q({open_n64320,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjax6 }));  // ../RTL/cortexm0ds_logic.v(18647)
  // ../RTL/cortexm0ds_logic.v(17815)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~B*~(D*A))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111001111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6684|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6_reg  (
    .a({open_n64321,_al_u5053_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u6683_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 ,_al_u6684_o}),
    .clk(XTAL1_wire),
    .d({_al_u5049_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dpwpw6 }),
    .f({_al_u6684_o,open_n64336}),
    .q({open_n64340,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 }));  // ../RTL/cortexm0ds_logic.v(17815)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u6688|_al_u6686  (
    .a({_al_u6686_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .b({_al_u6687_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hf0bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxrpw6 }),
    .f({_al_u6688_o,_al_u6686_o}));
  // ../RTL/cortexm0ds_logic.v(19125)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6693|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6_reg  (
    .a({_al_u6689_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 }),
    .b({_al_u6690_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 }),
    .c({_al_u6691_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6692_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 }),
    .mi({open_n64371,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6693_o,_al_u6691_o}),
    .q({open_n64375,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmzax6 }));  // ../RTL/cortexm0ds_logic.v(19125)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6694|_al_u6718  (
    .a({_al_u6688_o,_al_u6714_o}),
    .b({_al_u6693_o,_al_u6717_o}),
    .c({_al_u5031_o,_al_u5031_o}),
    .d({_al_u5260_o,_al_u5260_o}),
    .f({_al_u6694_o,_al_u6718_o}));
  // ../RTL/cortexm0ds_logic.v(18087)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6697|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 ,open_n64400}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4138_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 ,_al_u4136_o}),
    .f({_al_u6697_o,open_n64415}),
    .q({open_n64419,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z47ax6 }));  // ../RTL/cortexm0ds_logic.v(18087)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("(C*A*~(D*B))"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("(C*A*~(D*B))"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0010000010100000),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6698|_al_u7143  (
    .a({_al_u6696_o,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,_al_u4290_o}),
    .c({_al_u6697_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [14]}),
    .f({_al_u6698_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idkow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(C*B*~(D*~A))"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(C*B*~(D*~A))"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b1000000011000000),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b1000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6701|_al_u6700  (
    .a({_al_u4906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 }),
    .b({_al_u6698_o,_al_u6699_o}),
    .c({_al_u6700_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Heaax6 }),
    .f({_al_u6701_o,_al_u6700_o}));
  // ../RTL/cortexm0ds_logic.v(18088)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~B*~(D*A))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111001111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6703|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6_reg  (
    .a({open_n64468,_al_u5053_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u6702_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 ,_al_u6703_o}),
    .clk(XTAL1_wire),
    .d({_al_u5050_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ad7ax6 }),
    .f({_al_u6703_o,open_n64483}),
    .q({open_n64487,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 }));  // ../RTL/cortexm0ds_logic.v(18088)
  // ../RTL/cortexm0ds_logic.v(18577)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~D*~(~C*~A)))"),
    //.LUTF1("(~D*~(B*~(~C*~A)))"),
    //.LUTG0("(~B*~(~D*~(~C*~A)))"),
    //.LUTG1("(~D*~(B*~(~C*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100000001),
    .INIT_LUTF1(16'b0000000000110111),
    .INIT_LUTG0(16'b0011001100000001),
    .INIT_LUTG1(16'b0000000000110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6706|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 ,_al_u6596_o}),
    .b({_al_u1299_o,_al_u6706_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6706_o,open_n64505}),
    .q({open_n64509,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bciax6 }));  // ../RTL/cortexm0ds_logic.v(18577)
  // ../RTL/cortexm0ds_logic.v(18121)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6708|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u1699_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u5050_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .f({_al_u6708_o,open_n64530}),
    .q({open_n64534,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 }));  // ../RTL/cortexm0ds_logic.v(18121)
  // ../RTL/cortexm0ds_logic.v(18120)
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(C*~(D*B)))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(A*~(C*~(D*B)))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111010111110101),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0111010111110101),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6709|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6_reg  (
    .a({open_n64535,_al_u6709_o}),
    .b({_al_u6708_o,_al_u6719_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvabx6 ,_al_u5020_o}),
    .clk(XTAL1_wire),
    .d({_al_u5053_o,_al_u6725_o}),
    .f({_al_u6709_o,open_n64554}),
    .q({open_n64558,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sd8ax6 }));  // ../RTL/cortexm0ds_logic.v(18120)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6711|_al_u6710  (
    .a({open_n64559,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 }),
    .d({_al_u6710_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 }),
    .f({_al_u6711_o,_al_u6710_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6714|_al_u6712  (
    .a({open_n64584,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 }),
    .b({_al_u6712_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .c({_al_u6713_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K94bx6 }),
    .d({_al_u6711_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdxax6 }),
    .f({_al_u6714_o,_al_u6712_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u6716|_al_u5265  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ohyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yqzax6 }),
    .f({_al_u6716_o,_al_u5265_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u6717|_al_u6715  (
    .a({_al_u6715_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .b({_al_u6716_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gd0bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J6zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xo1bx6 }),
    .f({_al_u6717_o,_al_u6715_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u6719|_al_u6946  (
    .b({_al_u6718_o,_al_u6945_o}),
    .c({_al_u5067_o,_al_u6819_o}),
    .d({_al_u6637_o,_al_u6719_o}),
    .f({_al_u6719_o,_al_u6946_o}));
  // ../RTL/cortexm0ds_logic.v(19893)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*A*~(D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0010000010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6722|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6_reg  (
    .a({_al_u6720_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .c({_al_u6721_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 }),
    .mi({open_n64677,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .f({_al_u6722_o,_al_u6721_o}),
    .q({open_n64682,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqabx6 }));  // ../RTL/cortexm0ds_logic.v(19893)
  // ../RTL/cortexm0ds_logic.v(19890)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6724|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvsiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({_al_u6723_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Buabx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sb8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 }),
    .mi({open_n64693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .f({_al_u6724_o,_al_u6723_o}),
    .q({open_n64698,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkabx6 }));  // ../RTL/cortexm0ds_logic.v(19890)
  // ../RTL/cortexm0ds_logic.v(18122)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6727|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u1697_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u5050_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .f({_al_u6727_o,open_n64715}),
    .q({open_n64719,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh8ax6 }));  // ../RTL/cortexm0ds_logic.v(18122)
  // ../RTL/cortexm0ds_logic.v(19888)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(C*~(D*B)))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111010111110101),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6728|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6_reg  (
    .a({open_n64720,_al_u6728_o}),
    .b({_al_u6727_o,_al_u6732_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 ,_al_u5020_o}),
    .clk(XTAL1_wire),
    .d({_al_u5053_o,_al_u6738_o}),
    .f({_al_u6728_o,open_n64735}),
    .q({open_n64739,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ggabx6 }));  // ../RTL/cortexm0ds_logic.v(19888)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6730|_al_u6729  (
    .a({open_n64740,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F0eow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7kpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fb0bx6 }),
    .d({_al_u6729_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rk1bx6 }),
    .f({_al_u6730_o,_al_u6729_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u6732|_al_u6731  (
    .b({_al_u6731_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({_al_u5067_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 }),
    .d({_al_u6649_o,_al_u6730_o}),
    .f({_al_u6732_o,_al_u6731_o}));
  // ../RTL/cortexm0ds_logic.v(18253)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*A*~(D*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*A*~(D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0010000010100000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6735|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6_reg  (
    .a({_al_u6733_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({_al_u6734_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpxax6 }),
    .mi({open_n64790,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .f({_al_u6735_o,_al_u6734_o}),
    .q({open_n64806,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4cax6 }));  // ../RTL/cortexm0ds_logic.v(18253)
  // ../RTL/cortexm0ds_logic.v(18167)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6737|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6_reg  (
    .a({_al_u6735_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1tiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ureax6 }),
    .mi({open_n64810,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .f({_al_u6737_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1tiu6 }),
    .q({open_n64826,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oi9ax6 }));  // ../RTL/cortexm0ds_logic.v(18167)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6741|_al_u6740  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6lax6 }),
    .c({_al_u6740_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u4169_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0iax6 }),
    .f({_al_u6741_o,_al_u6740_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6743|_al_u6742  (
    .c({_al_u6742_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .d({_al_u6628_o,_al_u6741_o}),
    .f({_al_u6743_o,_al_u6742_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u6746|_al_u6745  (
    .c({_al_u6741_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 }),
    .d({_al_u6745_o,_al_u6628_o}),
    .f({_al_u6746_o,_al_u6745_o}));
  // ../RTL/cortexm0ds_logic.v(17870)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~(D*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000011100001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6749|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R05iu6 ,open_n64905}),
    .b({_al_u4170_o,open_n64906}),
    .c({_al_u6741_o,_al_u6749_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 ,_al_u6745_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6749_o,open_n64920}),
    .q({open_n64924,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7ypw6 }));  // ../RTL/cortexm0ds_logic.v(17870)
  // ../RTL/cortexm0ds_logic.v(19758)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6751|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 ,open_n64925}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 ,_al_u4052_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jl8iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F2dax6 ,_al_u4035_o}),
    .f({_al_u6751_o,open_n64944}),
    .q({open_n64948,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dm6bx6 }));  // ../RTL/cortexm0ds_logic.v(19758)
  // ../RTL/cortexm0ds_logic.v(18254)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*A*~(D*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*A*~(D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0010000010100000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6753|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6_reg  (
    .a({_al_u6751_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .c({_al_u6752_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Biaax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 }),
    .mi({open_n64952,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .f({_al_u6753_o,_al_u6752_o}),
    .q({open_n64968,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6cax6 }));  // ../RTL/cortexm0ds_logic.v(18254)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*~C*B))"),
    //.LUT1("(C*B*~(D*~A))"),
    .INIT_LUT0(16'b1010101010100010),
    .INIT_LUT1(16'b1000000011000000),
    .MODE("LOGIC"))
    \_al_u6756|_al_u5046  (
    .a({_al_u4816_o,_al_u5044_o}),
    .b({_al_u6755_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mmqiu6 }),
    .c({_al_u5044_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di3qw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Le2qw6 }),
    .f({_al_u6756_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }));
  // ../RTL/cortexm0ds_logic.v(17226)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~A*~(~C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110101110),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6758|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,_al_u2077_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 ,_al_u1892_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 ,_al_u2084_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 ,_al_u2085_o}),
    .f({_al_u6758_o,\u_cmsdk_mcu/HWDATA [12]}),
    .q({open_n65005,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyipw6 }));  // ../RTL/cortexm0ds_logic.v(17226)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~(D*A)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*~(C*~(D*A)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b1000110000001100),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1000110000001100),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6759|_al_u6913  (
    .a({_al_u6757_o,_al_u6626_o}),
    .b({_al_u6758_o,_al_u6819_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M0eow6 ,_al_u6759_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z71bx6 ,_al_u5067_o}),
    .f({_al_u6759_o,_al_u6913_o}));
  // ../RTL/cortexm0ds_logic.v(18131)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*B*~(D*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*B*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0100000011000000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6760|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6_reg  (
    .a({_al_u6626_o,open_n65030}),
    .b({_al_u6756_o,_al_u6762_o}),
    .c({_al_u6759_o,_al_u5020_o}),
    .clk(XTAL1_wire),
    .d({_al_u5067_o,_al_u6760_o}),
    .f({_al_u6760_o,open_n65049}),
    .q({open_n65053,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 }));  // ../RTL/cortexm0ds_logic.v(18131)
  // ../RTL/cortexm0ds_logic.v(18134)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6761|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,_al_u6761_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({_al_u5050_o,_al_u5053_o}),
    .mi({open_n65066,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .f({_al_u6761_o,_al_u6762_o}),
    .q({open_n65071,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Su8ax6 }));  // ../RTL/cortexm0ds_logic.v(18134)
  // ../RTL/cortexm0ds_logic.v(17412)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(~C*D))"),
    //.LUTF1("(~(D*~C)*~(B)*~(A)+~(D*~C)*B*~(A)+~(~(D*~C))*B*A+~(D*~C)*B*A)"),
    //.LUTG0("~(B*~(~C*D))"),
    //.LUTG1("(~(D*~C)*~(B)*~(A)+~(D*~C)*B*~(A)+~(~(D*~C))*B*A+~(D*~C)*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100110011),
    .INIT_LUTF1(16'b1101100011011101),
    .INIT_LUTG0(16'b0011111100110011),
    .INIT_LUTG1(16'b1101100011011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6765|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6_reg  (
    .a({_al_u6628_o,open_n65072}),
    .b({_al_u6649_o,_al_u6765_o}),
    .c({_al_u6742_o,_al_u4581_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ,_al_u6744_o}),
    .f({_al_u6765_o,open_n65091}),
    .q({open_n65095,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 }));  // ../RTL/cortexm0ds_logic.v(17412)
  // ../RTL/cortexm0ds_logic.v(17437)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(~C*D))"),
    //.LUTF1("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    //.LUTG0("~(B*~(~C*D))"),
    //.LUTG1("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100110011),
    .INIT_LUTF1(16'b0111001001110111),
    .INIT_LUTG0(16'b0011111100110011),
    .INIT_LUTG1(16'b0111001001110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6767|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6_reg  (
    .a({_al_u6628_o,open_n65096}),
    .b({_al_u6637_o,_al_u6767_o}),
    .c({_al_u6742_o,_al_u4611_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ,_al_u6744_o}),
    .f({_al_u6767_o,open_n65115}),
    .q({open_n65119,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 }));  // ../RTL/cortexm0ds_logic.v(17437)
  // ../RTL/cortexm0ds_logic.v(17208)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(~C*D))"),
    //.LUT1("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100110011),
    .INIT_LUT1(16'b0111001001110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6769|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6_reg  (
    .a({_al_u6628_o,open_n65120}),
    .b({_al_u6633_o,_al_u6769_o}),
    .c({_al_u6742_o,_al_u4637_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ,_al_u6744_o}),
    .f({_al_u6769_o,open_n65135}),
    .q({open_n65139,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 }));  // ../RTL/cortexm0ds_logic.v(17208)
  // ../RTL/cortexm0ds_logic.v(18563)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(~C*D))"),
    //.LUTF1("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    //.LUTG0("~(B*~(~C*D))"),
    //.LUTG1("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100110011),
    .INIT_LUTF1(16'b0111001001110111),
    .INIT_LUTG0(16'b0011111100110011),
    .INIT_LUTG1(16'b0111001001110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6771|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6_reg  (
    .a({_al_u6628_o,open_n65140}),
    .b({_al_u6650_o,_al_u6771_o}),
    .c({_al_u6742_o,_al_u4663_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ,_al_u6744_o}),
    .f({_al_u6771_o,open_n65159}),
    .q({open_n65163,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 }));  // ../RTL/cortexm0ds_logic.v(18563)
  // ../RTL/cortexm0ds_logic.v(18564)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(~C*D))"),
    //.LUT1("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100110011),
    .INIT_LUT1(16'b0111001001110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6773|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6_reg  (
    .a({_al_u6628_o,open_n65164}),
    .b({_al_u6652_o,_al_u6773_o}),
    .c({_al_u6742_o,_al_u4688_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ,_al_u6744_o}),
    .f({_al_u6773_o,open_n65179}),
    .q({open_n65183,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 }));  // ../RTL/cortexm0ds_logic.v(18564)
  // ../RTL/cortexm0ds_logic.v(18566)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b0011000111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6776|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6_reg  (
    .a({_al_u6744_o,open_n65184}),
    .b({_al_u6746_o,_al_u6776_o}),
    .c({_al_u4712_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [1]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 ,_al_u6775_o}),
    .f({_al_u6776_o,open_n65199}),
    .q({open_n65203,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8iax6 }));  // ../RTL/cortexm0ds_logic.v(18566)
  // ../RTL/cortexm0ds_logic.v(18621)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b0011000111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6778|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6_reg  (
    .a({_al_u6744_o,open_n65204}),
    .b({_al_u6746_o,_al_u6778_o}),
    .c({_al_u4735_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [2]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 ,_al_u6775_o}),
    .f({_al_u6778_o,open_n65219}),
    .q({open_n65223,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zqiax6 }));  // ../RTL/cortexm0ds_logic.v(18621)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u677|_al_u676  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vygax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .f({_al_u677_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I6row6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(18622)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("(~(D*B)*~(~C*A))"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b0011000111110101),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b0011000111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6780|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6_reg  (
    .a({_al_u6744_o,open_n65252}),
    .b({_al_u6746_o,_al_u6780_o}),
    .c({_al_u4836_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [3]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 ,_al_u6775_o}),
    .f({_al_u6780_o,open_n65271}),
    .q({open_n65275,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ysiax6 }));  // ../RTL/cortexm0ds_logic.v(18622)
  // ../RTL/cortexm0ds_logic.v(18623)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("(~(D*B)*~(~C*A))"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b0011000111110101),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b0011000111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6782|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6_reg  (
    .a({_al_u6744_o,open_n65276}),
    .b({_al_u6746_o,_al_u6782_o}),
    .c({_al_u4756_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [4]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 ,_al_u6775_o}),
    .f({_al_u6782_o,open_n65295}),
    .q({open_n65299,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuiax6 }));  // ../RTL/cortexm0ds_logic.v(18623)
  // ../RTL/cortexm0ds_logic.v(18624)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b0011000111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6784|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6_reg  (
    .a({_al_u6744_o,open_n65300}),
    .b({_al_u6746_o,_al_u6784_o}),
    .c({_al_u4776_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [5]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 ,_al_u6775_o}),
    .f({_al_u6784_o,open_n65315}),
    .q({open_n65319,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wwiax6 }));  // ../RTL/cortexm0ds_logic.v(18624)
  // ../RTL/cortexm0ds_logic.v(18625)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b0011000111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6786|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6_reg  (
    .a({_al_u6744_o,open_n65320}),
    .b({_al_u6746_o,_al_u6786_o}),
    .c({_al_u4796_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [6]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 ,_al_u6775_o}),
    .f({_al_u6786_o,open_n65335}),
    .q({open_n65339,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wyiax6 }));  // ../RTL/cortexm0ds_logic.v(18625)
  // ../RTL/cortexm0ds_logic.v(18626)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("(~(D*B)*~(~C*A))"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b0011000111110101),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b0011000111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6788|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6_reg  (
    .a({_al_u6744_o,open_n65340}),
    .b({_al_u6746_o,_al_u6788_o}),
    .c({_al_u4816_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [7]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 ,_al_u6775_o}),
    .f({_al_u6788_o,open_n65359}),
    .q({open_n65363,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0jax6 }));  // ../RTL/cortexm0ds_logic.v(18626)
  // ../RTL/cortexm0ds_logic.v(18627)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("(~(D*B)*~(~C*A))"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b0011000111110101),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b0011000111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6790|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6_reg  (
    .a({_al_u6744_o,open_n65364}),
    .b({_al_u6746_o,_al_u6790_o}),
    .c({_al_u4886_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [8]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 ,_al_u6775_o}),
    .f({_al_u6790_o,open_n65383}),
    .q({open_n65387,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W2jax6 }));  // ../RTL/cortexm0ds_logic.v(18627)
  // ../RTL/cortexm0ds_logic.v(17650)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(~C*D))"),
    //.LUT1("~((D*~C)*~(B)*~(A)+(D*~C)*B*~(A)+~((D*~C))*B*A+(D*~C)*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100110011),
    .INIT_LUT1(16'b0111001001110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6792|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6_reg  (
    .a({_al_u6628_o,open_n65388}),
    .b({_al_u6626_o,_al_u6792_o}),
    .c({_al_u6742_o,_al_u4865_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ,_al_u6744_o}),
    .f({_al_u6792_o,open_n65403}),
    .q({open_n65407,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 }));  // ../RTL/cortexm0ds_logic.v(17650)
  // ../RTL/cortexm0ds_logic.v(19970)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6794|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6_reg  (
    .a({_al_u5053_o,open_n65408}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sf1iu6 ,open_n65409}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 ,_al_u6812_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ,_al_u6794_o}),
    .f({_al_u6794_o,open_n65428}),
    .q({open_n65432,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8dbx6 }));  // ../RTL/cortexm0ds_logic.v(19970)
  // ../RTL/cortexm0ds_logic.v(18685)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    //.LUT1("(~(D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110100000001),
    .INIT_LUT1(16'b0011000111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6796|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wz4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iv1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qqhiu6 }),
    .c({_al_u1848_o,_al_u1848_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 }),
    .f({_al_u6796_o,open_n65447}),
    .q({open_n65451,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O2kax6 }));  // ../RTL/cortexm0ds_logic.v(18685)
  // ../RTL/cortexm0ds_logic.v(20099)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6801|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6_reg  (
    .a({_al_u6796_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .b({_al_u6798_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({_al_u6799_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6800_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 }),
    .mi({open_n65462,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .f({_al_u6801_o,_al_u6800_o}),
    .q({open_n65467,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzgbx6 }));  // ../RTL/cortexm0ds_logic.v(20099)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C*~B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(A*~(D*C*~B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1000101010101010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1000101010101010),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6802|_al_u6812  (
    .a({open_n65468,_al_u5020_o}),
    .b({open_n65469,_al_u6795_o}),
    .c({_al_u6801_o,_al_u6802_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 ,_al_u6811_o}),
    .f({_al_u6802_o,_al_u6812_o}));
  // ../RTL/cortexm0ds_logic.v(19617)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6805|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6_reg  (
    .a({_al_u6803_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smnow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K65bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 }),
    .mi({open_n65497,\u_cmsdk_mcu/HWDATA [23]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6805_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Smnow6 }),
    .q({open_n65512,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Od4bx6 }));  // ../RTL/cortexm0ds_logic.v(19617)
  // ../RTL/cortexm0ds_logic.v(19119)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6808|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6_reg  (
    .a({open_n65513,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 }),
    .b({_al_u6806_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvgiu6 }),
    .c({_al_u6807_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6805_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 }),
    .mi({open_n65524,\u_cmsdk_mcu/HWDATA [23]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6808_o,_al_u6807_o}),
    .q({open_n65528,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkzax6 }));  // ../RTL/cortexm0ds_logic.v(19119)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6809|_al_u2312  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8eiu6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L9eiu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J7xax6 }),
    .f({_al_u6809_o,_al_u2312_o}));
  // ../RTL/cortexm0ds_logic.v(18583)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(D*C*B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(~A*~(D*C*B))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110101010101010),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1110101010101010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u680|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6_reg  (
    .a({_al_u677_o,_al_u680_o}),
    .b({_al_u678_o,_al_u681_o}),
    .c({_al_u679_o,_al_u682_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u680_o,open_n65569}),
    .q({open_n65573,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdiax6 }));  // ../RTL/cortexm0ds_logic.v(18583)
  // ../RTL/cortexm0ds_logic.v(19017)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u6811|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6_reg  (
    .a({open_n65574,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 }),
    .b({_al_u6809_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 }),
    .c({_al_u6810_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nazax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6808_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 }),
    .mi({open_n65585,\u_cmsdk_mcu/HWDATA [23]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6811_o,_al_u6810_o}),
    .q({open_n65589,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slyax6 }));  // ../RTL/cortexm0ds_logic.v(19017)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*D))"),
    //.LUTF1("(D*~(C*~B*~A))"),
    //.LUTG0("(~C*~(B*D))"),
    //.LUTG1("(D*~(C*~B*~A))"),
    .INIT_LUTF0(16'b0000001100001111),
    .INIT_LUTF1(16'b1110111100000000),
    .INIT_LUTG0(16'b0000001100001111),
    .INIT_LUTG1(16'b1110111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6815|_al_u6814  (
    .a({_al_u677_o,open_n65590}),
    .b({_al_u3115_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv }),
    .c({_al_u6814_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P5vpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpnpw6 ,_al_u1658_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ,_al_u6814_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6816|_al_u6819  (
    .c({_al_u5001_o,_al_u5001_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ,_al_u6819_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(B*~(D*~(C*~A)))"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b0100000011001100),
    .MODE("LOGIC"))
    \_al_u6820|_al_u6818  (
    .a({_al_u6795_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha3ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjnow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .c({_al_u6811_o,_al_u6817_o}),
    .d({_al_u6819_o,_al_u1848_o}),
    .f({_al_u6820_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjnow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*C)*~(B*~A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b1011101100001011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u6822|_al_u6821  (
    .a({open_n65659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rw1iu6 }),
    .b({_al_u6821_o,_al_u6819_o}),
    .c({_al_u6817_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mg3ju6_lutinv ,_al_u1865_o}),
    .f({_al_u6822_o,_al_u6821_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~B)*~(A)*~(D)+(C*~B)*A*~(D)+~((C*~B))*A*D+(C*~B)*A*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~((C*~B)*~(A)*~(D)+(C*~B)*A*~(D)+~((C*~B))*A*D+(C*~B)*A*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0101010111001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0101010111001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6824|_al_u6823  (
    .a({open_n65680,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv }),
    .b({open_n65681,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({_al_u6823_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 }),
    .d({_al_u6822_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u6824_o,_al_u6823_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6825|_al_u4042  (
    .b({open_n65708,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0jiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owoiu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 }),
    .f({_al_u6825_o,_al_u4042_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*~C))"),
    //.LUT1("(D*~(~B*~(C*~A)))"),
    .INIT_LUT0(16'b0100010001000000),
    .INIT_LUT1(16'b1101110000000000),
    .MODE("LOGIC"))
    \_al_u6826|_al_u7053  (
    .a({_al_u6820_o,_al_u7013_o}),
    .b({_al_u6824_o,_al_u7052_o}),
    .c({_al_u6825_o,_al_u6820_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 }),
    .f({_al_u6826_o,_al_u7053_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6827|_al_u6702  (
    .b({open_n65755,_al_u6695_o}),
    .c({_al_u6819_o,_al_u6701_o}),
    .d({_al_u6695_o,_al_u5020_o}),
    .f({_al_u6827_o,_al_u6702_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D*~A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*~B)*~(D*~A))"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b1000101011001111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b1000101011001111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6829|_al_u6828  (
    .a({open_n65776,_al_u4735_o}),
    .b({_al_u6828_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxriu6 }),
    .c({_al_u6817_o,_al_u6819_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jb3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u6829_o,_al_u6828_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6831|_al_u7015  (
    .b({open_n65803,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv ,_al_u7015_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    //.LUT1("(~C*~B*~(~D*~A))"),
    .INIT_LUT0(16'b0000110011011101),
    .INIT_LUT1(16'b0000001100000010),
    .MODE("LOGIC"))
    \_al_u6833|_al_u6832  (
    .a({_al_u6829_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qdhow6_lutinv }),
    .b({_al_u6021_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({_al_u6830_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u6832_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u6833_o,_al_u6832_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(~C*~A))"),
    //.LUT1("(B*~(~D*~(C*~A)))"),
    .INIT_LUT0(16'b0011001011111010),
    .INIT_LUT1(16'b1100110001000000),
    .MODE("LOGIC"))
    \_al_u6836|_al_u6835  (
    .a({_al_u6827_o,_al_u6823_o}),
    .b({_al_u6833_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2ziu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bimow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u6836_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bimow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6838|_al_u698  (
    .b({_al_u698_o,open_n65866}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D31ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .d({_al_u1887_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u6838_o,_al_u698_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u6841|_al_u6840  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ,_al_u6219_o}),
    .f({_al_u6841_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6843|_al_u6842  (
    .c({_al_u6842_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .d({_al_u6841_o,_al_u6129_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxlow6 ,_al_u6842_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(D*C*~(B*~A))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b1011000000000000),
    .MODE("LOGIC"))
    \_al_u6844|_al_u7062  (
    .a({_al_u6826_o,open_n65943}),
    .b({_al_u6836_o,_al_u7060_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxlow6 ,_al_u6844_o}),
    .f({_al_u6844_o,_al_u7062_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*B)*~(D*A))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0101000111110011),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u6846|_al_u6845  (
    .a({open_n65964,_al_u6104_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .c({_al_u6819_o,_al_u1868_o}),
    .d({_al_u6676_o,_al_u6817_o}),
    .f({_al_u6846_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J9eow6 }));
  // ../RTL/cmsdk_apb_uart.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u684|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0],open_n65985}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [1],open_n65986}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3],_al_u685_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n40_lutinv ,open_n66003}),
    .q({open_n66007,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3]}));  // ../RTL/cmsdk_apb_uart.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D*~A))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~(C*~B)*~(D*~A))"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b1000101011001111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b1000101011001111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6851|_al_u6850  (
    .a({open_n66008,_al_u4836_o}),
    .b({_al_u6850_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4siu6 }),
    .c({_al_u6817_o,_al_u6819_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ,_al_u6850_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u6853|_al_u6852  (
    .a({open_n66033,_al_u4865_o}),
    .b({_al_u6852_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1xiu6 }),
    .c({_al_u6817_o,_al_u6819_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lj3ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u6853_o,_al_u6852_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0000010011000100),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0000010011000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6855|_al_u6932  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8viu6 ,_al_u1862_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U6wiu6 }),
    .c({_al_u5001_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv }),
    .d({_al_u1850_o,_al_u5001_o}),
    .f({_al_u6855_o,_al_u6932_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0000001111001111),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b0000001111001111),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6857|_al_u6976  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv }),
    .d({_al_u6129_o,_al_u6047_o}),
    .f({_al_u6857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*~A))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~(~D*B)*~(~C*~A))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111101000110010),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111101000110010),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6858|_al_u6854  (
    .a({open_n66104,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 }),
    .b({_al_u6856_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({_al_u6857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogdow6 ,_al_u6853_o}),
    .f({_al_u6858_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ogdow6 }));
  // ../RTL/cmsdk_apb_uart.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u685|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n40_lutinv ,open_n66131}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/baud_updated ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reload_i ,_al_u685_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u685_o,open_n66144}),
    .q({open_n66148,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [1]}));  // ../RTL/cmsdk_apb_uart.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6860|_al_u6859  (
    .a({open_n66149,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .b({open_n66150,_al_u2647_o}),
    .c({_al_u6859_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 }),
    .d({_al_u6841_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydopw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,_al_u6859_o}));
  // ../RTL/cortexm0ds_logic.v(18759)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~D)"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("~(C*B*~D)"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100111111),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6861|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Whmax6_reg  (
    .b({_al_u6858_o,_al_u6861_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdmiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6846_o,_al_u6844_o}),
    .f({_al_u6861_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .q({open_n66193,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[16] }));  // ../RTL/cortexm0ds_logic.v(18759)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6863|_al_u6865  (
    .c({_al_u6817_o,_al_u6817_o}),
    .d({_al_u5998_o,_al_u5998_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*C)*~(B*~A))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1011101100001011),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6866|_al_u6864  (
    .a({open_n66218,_al_u6057_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z4kow6 ,_al_u1833_o}),
    .f({_al_u6866_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z4kow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6867|_al_u6669  (
    .b({_al_u6866_o,_al_u6661_o}),
    .c({_al_u6819_o,_al_u6668_o}),
    .d({_al_u6661_o,_al_u5020_o}),
    .f({_al_u6867_o,_al_u6669_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(~A*~(C*B)))"),
    //.LUTG0("(~A*~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(~A*~(C*B)))"),
    .INIT_LUTF0(16'b0000010100010001),
    .INIT_LUTF1(16'b1110101000000000),
    .INIT_LUTG0(16'b0000010100010001),
    .INIT_LUTG1(16'b1110101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6868|_al_u6171  (
    .a({_al_u6171_o,_al_u6170_o}),
    .b({_al_u6170_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nweow6 }),
    .c({_al_u6021_o,_al_u6125_o}),
    .d({_al_u6817_o,_al_u5998_o}),
    .f({_al_u6868_o,_al_u6171_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b0000010011000100),
    .MODE("LOGIC"))
    \_al_u6869|_al_u5107  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 ,open_n66289}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfviu6 }),
    .c({_al_u5001_o,_al_u1852_o}),
    .d({_al_u1852_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u6869_o,_al_u5107_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(D*~(C*~B))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1100111100000000),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1100111100000000),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6872|_al_u6939  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ,_al_u6125_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv }),
    .d({_al_u6871_o,_al_u6938_o}),
    .f({_al_u6872_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6873|_al_u6955  (
    .b({_al_u6071_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .d({_al_u6872_o,_al_u6954_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D*~A))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(~(C*~B)*~(D*~A))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1000101011001111),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1000101011001111),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6875|_al_u6874  (
    .a({open_n66358,_al_u4581_o}),
    .b({_al_u6151_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovpiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,_al_u6819_o}),
    .d({_al_u6874_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u6875_o,_al_u6874_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(D*~(C*~B))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1100111100000000),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1100111100000000),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6876|_al_u6936  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ,_al_u6071_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv }),
    .d({_al_u6875_o,_al_u6935_o}),
    .f({_al_u6876_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*~A))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(~(~D*B)*~(~C*~A))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b1111101000110010),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111101000110010),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6878|_al_u6877  (
    .a({open_n66409,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bddow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({_al_u6857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 }),
    .d({_al_u6870_o,_al_u6876_o}),
    .f({_al_u6878_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bddow6 }));
  // ../RTL/cortexm0ds_logic.v(17708)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6879|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yhupw6_reg  (
    .b({_al_u6878_o,_al_u6879_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wamiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6867_o,_al_u6844_o}),
    .f({_al_u6879_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .q({open_n66452,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[15] }));  // ../RTL/cortexm0ds_logic.v(17708)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*D))"),
    //.LUTF1("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("(B*~(~C*D))"),
    //.LUTG1("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT_LUTF0(16'b1100000011001100),
    .INIT_LUTF1(16'b0000010011000100),
    .INIT_LUTG0(16'b1100000011001100),
    .INIT_LUTG1(16'b0000010011000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6882|_al_u5094  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 ,open_n66453}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wmviu6 }),
    .c({_al_u5001_o,_al_u1854_o}),
    .d({_al_u1854_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u6882_o,_al_u5094_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~A*~(C*B)))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(~A*~(C*B)))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1110101000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1110101000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6883|_al_u6881  (
    .a({open_n66478,_al_u6167_o}),
    .b({open_n66479,_al_u6166_o}),
    .c({_al_u6882_o,_al_u6021_o}),
    .d({_al_u6881_o,_al_u6817_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ,_al_u6881_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(C*~(D*~B)))"),
    //.LUTF1("(~(C*~B)*~(D*~A))"),
    //.LUTG0("(A*~(C*~(D*~B)))"),
    //.LUTG1("(~(C*~B)*~(D*~A))"),
    .INIT_LUTF0(16'b0010101000001010),
    .INIT_LUTF1(16'b1000101011001111),
    .INIT_LUTG0(16'b0010101000001010),
    .INIT_LUTG1(16'b1000101011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6884|_al_u5232  (
    .a({_al_u4776_o,_al_u5020_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bisiu6 ,_al_u4776_o}),
    .c({_al_u6819_o,_al_u5231_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({_al_u6884_o,_al_u5232_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6885|_al_u6919  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 ,_al_u6082_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv }),
    .d({_al_u6884_o,_al_u6918_o}),
    .f({_al_u6885_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(D*~(C*~B))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1100111100000000),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1100111100000000),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6886|_al_u6905  (
    .b({_al_u6068_o,_al_u6018_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .d({_al_u6885_o,_al_u6904_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6888|_al_u6887  (
    .a({open_n66576,_al_u4611_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 ,_al_u6819_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({_al_u6887_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jaqiu6 }),
    .f({_al_u6888_o,_al_u6887_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*C)*~(B*~A))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b1011101100001011),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u6892|_al_u6891  (
    .a({open_n66601,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U1uiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,_al_u6819_o}),
    .c({_al_u6891_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R04ju6 ,_al_u1836_o}),
    .f({_al_u6892_o,_al_u6891_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*~A))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1111101000110010),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u6894|_al_u6890  (
    .a({open_n66622,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 }),
    .b({_al_u6890_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 }),
    .f({_al_u6894_o,_al_u6890_o}));
  // ../RTL/cortexm0ds_logic.v(18757)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~D)"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("~(C*B*~D)"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100111111),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6895|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wdmax6_reg  (
    .b({_al_u6894_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 }),
    .c({_al_u6857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7miu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ,_al_u6844_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .q({open_n66665,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[18] }));  // ../RTL/cortexm0ds_logic.v(18757)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    //.LUT1("(D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b0001000100000101),
    .INIT_LUT1(16'b1110101000000000),
    .MODE("LOGIC"))
    \_al_u6897|_al_u6169  (
    .a({_al_u6169_o,_al_u6168_o}),
    .b({_al_u6168_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csnow6 }),
    .c({_al_u6021_o,_al_u6015_o}),
    .d({_al_u6817_o,_al_u5998_o}),
    .f({_al_u6897_o,_al_u6169_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000010011000100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6899|_al_u6898  (
    .a({open_n66686,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wtviu6 }),
    .b({open_n66687,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv }),
    .c({_al_u6898_o,_al_u5001_o}),
    .d({_al_u6897_o,_al_u1856_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ,_al_u6898_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6901|_al_u6900  (
    .a({open_n66708,_al_u4796_o}),
    .b({_al_u6064_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uosiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,_al_u6819_o}),
    .d({_al_u6900_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u6901_o,_al_u6900_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(D*~(C*~B))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1100111100000000),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1100111100000000),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6902|_al_u6909  (
    .b({_al_u6075_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C34ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv }),
    .d({_al_u6901_o,_al_u6908_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D*~A))"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~(C*~B)*~(D*~A))"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b1000101011001111),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b1000101011001111),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6904|_al_u6903  (
    .a({open_n66755,_al_u4637_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tmqiu6 }),
    .c({_al_u6903_o,_al_u6819_o}),
    .d({_al_u6139_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u6904_o,_al_u6903_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~(B*~D))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0000111100000011),
    .MODE("LOGIC"))
    \_al_u6908|_al_u6907  (
    .a({open_n66780,_al_u1839_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U8uiu6 }),
    .c({_al_u6907_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hemow6_lutinv }),
    .d({_al_u6086_o,_al_u5001_o}),
    .f({_al_u6908_o,_al_u6907_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*~A))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1111101000110010),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u6910|_al_u6906  (
    .a({open_n66801,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6dow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 }),
    .f({_al_u6910_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6dow6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~D))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~(~C*~D))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b1100110011000000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1100110011000000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6911|_al_u7113  (
    .b({_al_u6910_o,_al_u7112_o}),
    .c({_al_u6857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 ,_al_u7113_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*~A))"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~(~D*C)*~(B*~A))"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b1011101100001011),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6915|_al_u6914  (
    .a({open_n66848,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bguiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,_al_u6819_o}),
    .c({_al_u6914_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({_al_u6034_o,_al_u1841_o}),
    .f({_al_u6915_o,_al_u6914_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u6918|_al_u6917  (
    .a({open_n66873,_al_u4663_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqiu6 }),
    .c({_al_u6917_o,_al_u6819_o}),
    .d({_al_u6135_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u6918_o,_al_u6917_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*C)*~(B*~A))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b1011101100001011),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u6922|_al_u6921  (
    .a({open_n66894,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0wiu6 }),
    .b({_al_u6921_o,_al_u6819_o}),
    .c({_al_u6817_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xa4ju6_lutinv ,_al_u1859_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ,_al_u6921_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*~A))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~(~D*B)*~(~C*~A))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111101000110010),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111101000110010),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6923|_al_u6920  (
    .a({open_n66915,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({_al_u6857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 }),
    .d({_al_u6920_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 }),
    .f({_al_u6923_o,_al_u6920_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(~D*~(C*~B))"),
    //.LUTG0("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(~D*~(C*~B))"),
    .INIT_LUTF0(16'b0011010100000000),
    .INIT_LUTF1(16'b0000000011001111),
    .INIT_LUTG0(16'b0011010100000000),
    .INIT_LUTG1(16'b0000000011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6925|_al_u6924  (
    .a({open_n66940,_al_u6061_o}),
    .b({_al_u4816_o,_al_u6079_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ,_al_u5998_o}),
    .d({_al_u6924_o,_al_u6817_o}),
    .f({_al_u6925_o,_al_u6924_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~(D*~A))"),
    //.LUT1("(~(D*~C)*~(B*~A))"),
    .INIT_LUT0(16'b1000000011000000),
    .INIT_LUT1(16'b1011000010111011),
    .MODE("LOGIC"))
    \_al_u6928|_al_u6738  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uc4ju6 ,_al_u4886_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yw1iu6 }),
    .c({_al_u4886_o,_al_u6737_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/St1iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxeow6 ,_al_u6738_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6929|_al_u6930  (
    .b({_al_u6057_o,_al_u6929_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,_al_u6819_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bxeow6 ,_al_u6732_o}),
    .f({_al_u6929_o,_al_u6930_o}));
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u692|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b0  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [0]}),
    .clk(1'b1),
    .d({_al_u566_o,_al_u3041_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u692_o,open_n67032}),
    .q({open_n67036,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [0]}));  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(C*B)))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1110101000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6933|_al_u6931  (
    .a({open_n67037,_al_u6163_o}),
    .b({open_n67038,_al_u6159_o}),
    .c({_al_u6932_o,_al_u6021_o}),
    .d({_al_u6931_o,_al_u6817_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ,_al_u6931_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6935|_al_u6934  (
    .a({open_n67059,_al_u4688_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mu3ju6 ,_al_u6819_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({_al_u6934_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eariu6 }),
    .f({_al_u6935_o,_al_u6934_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*~A))"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~(~D*C)*~(B*~A))"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b1011101100001011),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6938|_al_u6937  (
    .a({open_n67084,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Umuiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv ,_al_u6819_o}),
    .c({_al_u6937_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F14ju6 ,_al_u1844_o}),
    .f({_al_u6938_o,_al_u6937_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(~D*~A))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(~(~C*B)*~(~D*~A))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b1111001110100010),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111001110100010),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6941|_al_u6940  (
    .a({open_n67109,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nycow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({_al_u6857_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 }),
    .f({_al_u6941_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nycow6 }));
  // ../RTL/cortexm0ds_logic.v(18754)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(D*B*~(~C*~A))"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(D*B*~(~C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b1100100000000000),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b1100100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6942|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W7max6_reg  (
    .a({_al_u6930_o,open_n67134}),
    .b({_al_u6941_o,open_n67135}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ,_al_u6942_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Azliu6 ,_al_u6844_o}),
    .f({_al_u6942_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .q({open_n67156,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[21] }));  // ../RTL/cortexm0ds_logic.v(18754)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~C)*~(B*~A))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(~(D*~C)*~(B*~A))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b1011000010111011),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1011000010111011),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6945|_al_u6944  (
    .a({open_n67157,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Id4ju6 }),
    .b({_al_u6054_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,_al_u4529_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1low6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .f({_al_u6945_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1low6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*C)*~(B*~A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(~D*C)*~(B*~A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1011101100001011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1011101100001011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6949|_al_u6948  (
    .a({open_n67182,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bewiu6 }),
    .b({open_n67183,_al_u6819_o}),
    .c({_al_u6948_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({_al_u6947_o,_al_u1286_o}),
    .f({_al_u6949_o,_al_u6948_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u6951|_al_u6952  (
    .b({_al_u6068_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yt3ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qtfow6_lutinv }),
    .d({_al_u6950_o,_al_u6951_o}),
    .f({_al_u6951_o,_al_u6952_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*C)*~(B*~A))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b1011101100001011),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u6954|_al_u6953  (
    .a({open_n67230,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ntuiu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dyeow6_lutinv ,_al_u6819_o}),
    .c({_al_u6953_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q2eow6 }),
    .d({_al_u6122_o,_al_u1846_o}),
    .f({_al_u6954_o,_al_u6953_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*B)*~(~D*~A))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1111001110100010),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u6957|_al_u6956  (
    .a({open_n67251,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 }),
    .b({_al_u6956_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({_al_u6857_o,_al_u6952_o}),
    .d({_al_u6949_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 }),
    .f({_al_u6957_o,_al_u6956_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*~B))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(C*~A*~(~D*~B))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b0101000001000000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0101000001000000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6958|_al_u7049  (
    .a({open_n67272,_al_u7013_o}),
    .b({_al_u6957_o,_al_u6946_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ,_al_u7048_o}),
    .d({_al_u6946_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 }),
    .f({_al_u6958_o,_al_u7049_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0001001100110011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u695|_al_u2459  (
    .a({open_n67297,_al_u695_o}),
    .b({open_n67298,_al_u2458_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 ,_al_u1296_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .f({_al_u695_o,_al_u2459_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*~A))"),
    //.LUT1("(B*~(~C*~(D*~A)))"),
    .INIT_LUT0(16'b1111101000110010),
    .INIT_LUT1(16'b1100010011000000),
    .MODE("LOGIC"))
    \_al_u6961|_al_u6960  (
    .a({_al_u6827_o,_al_u6822_o}),
    .b({_al_u6960_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ,_al_u6857_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ,_al_u6829_o}),
    .f({_al_u6961_o,_al_u6960_o}));
  // ../RTL/cortexm0ds_logic.v(18970)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(D*~(~C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6962|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvxax6_reg  (
    .b({_al_u6820_o,_al_u6962_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evkiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6961_o,_al_u6844_o}),
    .f({_al_u6962_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .q({open_n67357,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] }));  // ../RTL/cortexm0ds_logic.v(18970)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~D))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~(~B*~D))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000011000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000011000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6964|_al_u2846  (
    .b({open_n67360,_al_u2845_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .d({_al_u6842_o,_al_u2843_o}),
    .f({_al_u6964_o,_al_u2846_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001111001111),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u6965|_al_u6847  (
    .b({_al_u6964_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .d({_al_u6047_o,_al_u6047_o}),
    .f({_al_u6965_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~B*~A*~(D*C))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000100010001),
    .MODE("LOGIC"))
    \_al_u6966|_al_u6243  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,open_n67407}),
    .b({_al_u6243_o,open_n67408}),
    .c({_al_u609_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .d({_al_u698_o,_al_u1662_o}),
    .f({_al_u6966_o,_al_u6243_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(~D*~C*B*~A)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(~D*~C*B*~A)"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b0000000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6967|_al_u6849  (
    .a({_al_u6841_o,open_n67429}),
    .b({_al_u6965_o,_al_u604_o}),
    .c({_al_u6848_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({_al_u6966_o,_al_u6848_o}),
    .f({_al_u6967_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~C*~(B*~D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0000111100000011),
    .MODE("LOGIC"))
    \_al_u6969|_al_u6968  (
    .b({_al_u6836_o,_al_u6830_o}),
    .c({_al_u6968_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .d({_al_u6826_o,_al_u6967_o}),
    .f({_al_u6969_o,_al_u6968_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6971|_al_u6970  (
    .c({_al_u1582_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u6970_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T23ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4mow6_lutinv ,_al_u6970_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*~(C)*D))"),
    //.LUT1("(A*~(~B*~(~D*C)))"),
    .INIT_LUT0(16'b0000000101000100),
    .INIT_LUT1(16'b1000100010101000),
    .MODE("LOGIC"))
    \_al_u6973|_al_u6972  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4mow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({_al_u6972_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,_al_u6972_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*~(~C*~A))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1111101011001000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u6978|_al_u6975  (
    .a({open_n67520,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 }),
    .b({_al_u6977_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 }),
    .d({_al_u6975_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 }),
    .f({_al_u6978_o,_al_u6975_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(B)*~((~C*A))*~(D)+~(B)*(~C*A)*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+B*(~C*A)*D)"),
    //.LUTF1("~((D*~C)*~(A)*~(B)+(D*~C)*A*~(B)+~((D*~C))*A*B+(D*~C)*A*B)"),
    //.LUTG0("(~(B)*~((~C*A))*~(D)+~(B)*(~C*A)*~(D)+~(B)*~((~C*A))*D+B*~((~C*A))*D+B*(~C*A)*D)"),
    //.LUTG1("~((D*~C)*~(A)*~(B)+(D*~C)*A*~(B)+~((D*~C))*A*B+(D*~C)*A*B)"),
    .INIT_LUTF0(16'b1111110100110011),
    .INIT_LUTF1(16'b0111010001110111),
    .INIT_LUTG0(16'b1111110100110011),
    .INIT_LUTG1(16'b0111010001110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6980|_al_u6979  (
    .a({_al_u6049_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .c({_al_u6979_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .f({_al_u6980_o,_al_u6979_o}));
  // ../RTL/cortexm0ds_logic.v(18763)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(D*~(~C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6981|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpmax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ,_al_u6981_o}),
    .c({_al_u6980_o,_al_u6183_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6978_o,_al_u6969_o}),
    .f({_al_u6981_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .q({open_n67583,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[10] }));  // ../RTL/cortexm0ds_logic.v(18763)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~B)*~(~C*~A))"),
    //.LUTF1("(C*~(~B*~(D*~A)))"),
    //.LUTG0("(~(~D*~B)*~(~C*~A))"),
    //.LUTG1("(C*~(~B*~(D*~A)))"),
    .INIT_LUTF0(16'b1111101011001000),
    .INIT_LUTF1(16'b1101000011000000),
    .INIT_LUTG0(16'b1111101011001000),
    .INIT_LUTG1(16'b1101000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6984|_al_u6983  (
    .a({_al_u6827_o,_al_u6822_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,_al_u6977_o}),
    .c({_al_u6983_o,_al_u6980_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ,_al_u6829_o}),
    .f({_al_u6984_o,_al_u6983_o}));
  // ../RTL/cortexm0ds_logic.v(19788)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~D)"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("~(C*B*~D)"),
    //.LUTG1("(D*~(~C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100111111),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6985|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zz7bx6_reg  (
    .b({_al_u6820_o,_al_u6985_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ngmiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6984_o,_al_u6969_o}),
    .f({_al_u6985_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .q({open_n67630,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[15] }));  // ../RTL/cortexm0ds_logic.v(19788)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(~D*~A))"),
    //.LUT1("(~(~D*~B)*~(~C*~A))"),
    .INIT_LUT0(16'b1111110010101000),
    .INIT_LUT1(16'b1111101011001000),
    .MODE("LOGIC"))
    \_al_u6987|_al_u7055  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,_al_u7016_o}),
    .b({_al_u6977_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 }),
    .d({_al_u6876_o,_al_u6876_o}),
    .f({_al_u6987_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt6ow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u6988|_al_u6994  (
    .b({_al_u6870_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 }),
    .c({_al_u6980_o,_al_u6980_o}),
    .d({_al_u6987_o,_al_u6993_o}),
    .f({_al_u6988_o,_al_u6994_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*~B))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(C*~A*~(~D*~B))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b0101000001000000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0101000001000000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6989|_al_u7105  (
    .a({open_n67673,_al_u7092_o}),
    .b({_al_u6988_o,_al_u6867_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ,_al_u7104_o}),
    .d({_al_u6867_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }),
    .f({_al_u6989_o,_al_u7105_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(~D*~A))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(~(~C*~B)*~(~D*~A))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b1111110010101000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111110010101000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6993|_al_u6992  (
    .a({open_n67698,_al_u6977_o}),
    .b({_al_u6992_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 }),
    .f({_al_u6993_o,_al_u6992_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~B)*~(~C*A))"),
    //.LUTF1("(~(~D*~B)*~(~C*~A))"),
    //.LUTG0("(~(~D*~B)*~(~C*A))"),
    //.LUTG1("(~(~D*~B)*~(~C*~A))"),
    .INIT_LUTF0(16'b1111010111000100),
    .INIT_LUTF1(16'b1111101011001000),
    .INIT_LUTG0(16'b1111010111000100),
    .INIT_LUTG1(16'b1111101011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6996|_al_u7099  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .b({_al_u6977_o,_al_u7093_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 }),
    .d({_al_u6853_o,_al_u6853_o}),
    .f({_al_u6996_o,_al_u7099_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6997|_al_u6856  (
    .b({_al_u6856_o,_al_u6855_o}),
    .c({_al_u6980_o,_al_u6817_o}),
    .d({_al_u6996_o,_al_u6036_o}),
    .f({_al_u6997_o,_al_u6856_o}));
  // ../RTL/cortexm0ds_logic.v(18765)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u6998|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtmax6_reg  (
    .b({_al_u6997_o,_al_u6998_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ,_al_u5918_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6846_o,_al_u6969_o}),
    .f({_al_u6998_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .q({open_n67791,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[8] }));  // ../RTL/cortexm0ds_logic.v(18765)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(~D*~A))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~(~C*~B)*~(~D*~A))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111110010101000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111110010101000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7001|_al_u7000  (
    .a({open_n67792,_al_u6977_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 }),
    .c({_al_u6980_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 }),
    .d({_al_u7000_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 }),
    .f({_al_u7001_o,_al_u7000_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~(D*~A)))"),
    //.LUTF1("(B*~(~C*~(D*~A)))"),
    //.LUTG0("(B*~(~C*~(D*~A)))"),
    //.LUTG1("(B*~(~C*~(D*~A)))"),
    .INIT_LUTF0(16'b1100010011000000),
    .INIT_LUTF1(16'b1100010011000000),
    .INIT_LUTG0(16'b1100010011000000),
    .INIT_LUTG1(16'b1100010011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7002|_al_u6926  (
    .a({_al_u6913_o,_al_u6913_o}),
    .b({_al_u7001_o,_al_u6923_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 }),
    .d({_al_u6925_o,_al_u6925_o}),
    .f({_al_u7002_o,_al_u6926_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~B)*~(~C*~A))"),
    //.LUTF1("(~(~D*~B)*~(~C*~A))"),
    //.LUTG0("(~(~D*~B)*~(~C*~A))"),
    //.LUTG1("(~(~D*~B)*~(~C*~A))"),
    .INIT_LUTF0(16'b1111101011001000),
    .INIT_LUTF1(16'b1111101011001000),
    .INIT_LUTG0(16'b1111101011001000),
    .INIT_LUTG1(16'b1111101011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7004|_al_u7043  (
    .a({_al_u6977_o,_al_u7016_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qodow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpeow6 }));
  // ../RTL/cortexm0ds_logic.v(18761)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~D)"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("~(C*B*~D)"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100111111),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u7006|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlmax6_reg  (
    .b({_al_u7005_o,_al_u7006_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,_al_u5954_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6930_o,_al_u6969_o}),
    .f({_al_u7006_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .q({open_n67887,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[13] }));  // ../RTL/cortexm0ds_logic.v(18761)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*~(~C*~A))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1111101011001000),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u7009|_al_u7008  (
    .a({open_n67888,_al_u6977_o}),
    .b({_al_u7008_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 }),
    .c({_al_u6980_o,_al_u6952_o}),
    .d({_al_u6949_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 }),
    .f({_al_u7009_o,_al_u7008_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u700|_al_u701  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Np7ow6_lutinv ,_al_u700_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae0iu6_lutinv }),
    .d({_al_u698_o,_al_u697_o}),
    .f({_al_u700_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u7010|_al_u7117  (
    .b({_al_u7009_o,_al_u7116_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkdow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .d({_al_u6946_o,_al_u6946_o}),
    .f({_al_u7010_o,_al_u7117_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("~(C*~((~B*~A))*~(D)+C*(~B*~A)*~(D)+~(C)*(~B*~A)*D+C*(~B*~A)*D)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("~(C*~((~B*~A))*~(D)+C*(~B*~A)*~(D)+~(C)*(~B*~A)*D+C*(~B*~A)*D)"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1110111000001111),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1110111000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7012|_al_u6047  (
    .a({_al_u6046_o,open_n67957}),
    .b({_al_u6100_o,_al_u604_o}),
    .c({_al_u6830_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,_al_u6046_o}),
    .f({_al_u7012_o,_al_u6047_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(D*B))"),
    //.LUTF1("(A*~(~B*~(~D*C)))"),
    //.LUTG0("(C*~A*~(D*B))"),
    //.LUTG1("(A*~(~B*~(~D*C)))"),
    .INIT_LUTF0(16'b0001000001010000),
    .INIT_LUTF1(16'b1000100010101000),
    .INIT_LUTG0(16'b0001000001010000),
    .INIT_LUTG1(16'b1000100010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7016|_al_u7014  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eccow6 ,_al_u6970_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aujpw6 }),
    .c({_al_u7014_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3vpw6 }),
    .d({_al_u7015_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzupw6 }),
    .f({_al_u7016_o,_al_u7014_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C*~B))"),
    //.LUTF1("(~A*~(~B*~(D*C)))"),
    //.LUTG0("(A*~(D*C*~B))"),
    //.LUTG1("(~A*~(~B*~(D*C)))"),
    .INIT_LUTF0(16'b1000101010101010),
    .INIT_LUTF1(16'b0101010001000100),
    .INIT_LUTG0(16'b1000101010101010),
    .INIT_LUTG1(16'b0101010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7018|_al_u6977  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .c({_al_u1658_o,_al_u1658_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pthiu6 }),
    .f({_al_u7018_o,_al_u6977_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~A*~(~D*B))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~A*~(~D*B))"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010100000001),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7019|_al_u6974  (
    .a({_al_u6964_o,open_n68030}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .c({_al_u7018_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ,_al_u6964_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kldow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0001000000010011),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u7021|_al_u7022  (
    .a({open_n68055,_al_u6046_o}),
    .b({open_n68056,_al_u7021_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .f({_al_u7021_o,_al_u7022_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(~D*~A))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1111110010101000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u7023|_al_u7020  (
    .a({open_n68077,_al_u7016_o}),
    .b({_al_u6856_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 }),
    .c({_al_u7022_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rcliu6 }),
    .d({_al_u7020_o,_al_u6853_o}),
    .f({_al_u7023_o,_al_u7020_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(~(~D*B)*~(C*A))"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(~(~D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b0101111100010011),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b0101111100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7024|_al_u7017  (
    .a({_al_u1658_o,open_n68098}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbhow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldiow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S4kbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .f({_al_u7024_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G8how6 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(~C*~(~B*D))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(~C*~(~B*D))"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b0000110000001111),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b0000110000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7026|_al_u7025  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R3how6_lutinv ,_al_u7024_o}),
    .c({_al_u7025_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ms5bx6 }),
    .d({_al_u6848_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ,_al_u7025_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7028|_al_u7013  (
    .b({open_n68151,_al_u6836_o}),
    .c({_al_u7027_o,_al_u7012_o}),
    .d({_al_u7013_o,_al_u6826_o}),
    .f({_al_u7028_o,_al_u7013_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0011000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u702|_al_u1314  (
    .b({open_n68178,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,_al_u702_o}),
    .f({_al_u702_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(~D*~A))"),
    //.LUTF1("(~(~C*~B)*~(~D*~A))"),
    //.LUTG0("(~(~C*~B)*~(~D*~A))"),
    //.LUTG1("(~(~C*~B)*~(~D*~A))"),
    .INIT_LUTF0(16'b1111110010101000),
    .INIT_LUTF1(16'b1111110010101000),
    .INIT_LUTG0(16'b1111110010101000),
    .INIT_LUTG1(16'b1111110010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7030|_al_u7034  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 }),
    .f({_al_u7030_o,_al_u7034_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(~D*~C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(~D*~C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b0100010001000000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0100010001000000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7031|_al_u7032  (
    .a({open_n68223,_al_u7013_o}),
    .b({_al_u7030_o,_al_u7031_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 }),
    .d({_al_u7016_o,_al_u7022_o}),
    .f({_al_u7031_o,_al_u7032_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*~C))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b0100010001000000),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u7035|_al_u7036  (
    .a({open_n68248,_al_u7013_o}),
    .b({_al_u7034_o,_al_u7035_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfcow6 }),
    .d({_al_u7016_o,_al_u7022_o}),
    .f({_al_u7035_o,_al_u7036_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(~D*~A))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1111110010101000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u7039|_al_u7038  (
    .a({open_n68269,_al_u7016_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 }),
    .c({_al_u7022_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 }),
    .d({_al_u7038_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 }),
    .f({_al_u7039_o,_al_u7038_o}));
  // ../RTL/cortexm0ds_logic.v(18713)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u703|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2lax6_reg  (
    .a({open_n68290,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u702_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[0] }),
    .mi({open_n68301,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,_al_u705_o}),
    .q({open_n68306,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[0] }));  // ../RTL/cortexm0ds_logic.v(18713)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~(D*~A)))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(~C*~(D*~A)))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1100010011000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100010011000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7041|_al_u7040  (
    .a({open_n68307,_al_u6913_o}),
    .b({open_n68308,_al_u7039_o}),
    .c({_al_u7040_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 }),
    .d({_al_u7013_o,_al_u6925_o}),
    .f({_al_u7041_o,_al_u7040_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*~B))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(C*~A*~(~D*~B))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0101000001000000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0101000001000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7044|_al_u7045  (
    .a({open_n68333,_al_u7013_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ,_al_u6930_o}),
    .c({_al_u7022_o,_al_u7044_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpeow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 }),
    .f({_al_u7044_o,_al_u7045_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~B)*~(~C*~A))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(~(~D*~B)*~(~C*~A))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b1111101011001000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111101011001000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7048|_al_u7047  (
    .a({open_n68358,_al_u7016_o}),
    .b({_al_u7047_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 }),
    .c({_al_u7022_o,_al_u6952_o}),
    .d({_al_u6949_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 }),
    .f({_al_u7048_o,_al_u7047_o}));
  // ../RTL/cortexm0ds_logic.v(17552)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u704|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9qpw6_reg  (
    .a({open_n68383,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u702_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] }),
    .mi({open_n68387,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ,_al_u819_o}),
    .q({open_n68403,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[28] }));  // ../RTL/cortexm0ds_logic.v(17552)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(~D*~A))"),
    //.LUTF1("(B*~(~C*~(D*~A)))"),
    //.LUTG0("(~(~C*~B)*~(~D*~A))"),
    //.LUTG1("(B*~(~C*~(D*~A)))"),
    .INIT_LUTF0(16'b1111110010101000),
    .INIT_LUTF1(16'b1100010011000000),
    .INIT_LUTG0(16'b1111110010101000),
    .INIT_LUTG1(16'b1100010011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7052|_al_u7051  (
    .a({_al_u6827_o,_al_u7016_o}),
    .b({_al_u7051_o,_al_u6822_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ycliu6 ,_al_u7022_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 ,_al_u6829_o}),
    .f({_al_u7052_o,_al_u7051_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*~B))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(C*~A*~(~D*~B))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0101000001000000),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0101000001000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7056|_al_u7057  (
    .a({open_n68428,_al_u7013_o}),
    .b({_al_u6870_o,_al_u6867_o}),
    .c({_al_u7022_o,_al_u7056_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mt6ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfliu6 }),
    .f({_al_u7056_o,_al_u7057_o}));
  // ../RTL/cortexm0ds_logic.v(18736)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111001101010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0111001101010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7059|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6_reg  (
    .a({_al_u1774_o,_al_u1796_o}),
    .b({_al_u1791_o,_al_u1794_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 ,_al_u1797_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qakbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7059_o,open_n68470}),
    .q({open_n68474,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Halax6 }));  // ../RTL/cortexm0ds_logic.v(18736)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTF1("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUTG1("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT_LUTF0(16'b0010011110101111),
    .INIT_LUTF1(16'b0010011110101111),
    .INIT_LUTG0(16'b0010011110101111),
    .INIT_LUTG1(16'b0010011110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7064|_al_u7189  (
    .a({_al_u4289_o,_al_u4289_o}),
    .b({_al_u4290_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [21],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [12]}),
    .f({_al_u7064_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hndow6 }));
  // ../RTL/cortexm0ds_logic.v(19901)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*A*~(D*~B))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111101011111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7065|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxabx6_reg  (
    .a({open_n68499,_al_u7062_o}),
    .b({_al_u7064_o,_al_u6958_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23],_al_u7065_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7065_o,open_n68513}),
    .q({open_n68517,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] }));  // ../RTL/cortexm0ds_logic.v(19901)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u7067|_al_u7186  (
    .a({open_n68518,_al_u4289_o}),
    .b({open_n68519,_al_u4290_o}),
    .c({_al_u4290_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] }),
    .d({_al_u4289_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [11]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Prdow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0010011110101111),
    .MODE("LOGIC"))
    \_al_u7068|_al_u7063  (
    .a({_al_u4289_o,open_n68540}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ,open_n68541}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17],_al_u4289_o}),
    .f({_al_u7068_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 }));
  // ../RTL/cortexm0ds_logic.v(18501)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*A*~(D*~B))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111101011111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7069|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thhax6_reg  (
    .a({open_n68562,_al_u7062_o}),
    .b({_al_u7068_o,_al_u6861_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [15],_al_u7069_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7069_o,open_n68576}),
    .q({open_n68580,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] }));  // ../RTL/cortexm0ds_logic.v(18501)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0010011110101111),
    .MODE("LOGIC"))
    \_al_u7071|_al_u7074  (
    .a({_al_u4289_o,_al_u4289_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19]}),
    .f({_al_u7071_o,_al_u7074_o}));
  // ../RTL/cortexm0ds_logic.v(18495)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*A*~(D*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(C*A*~(D*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0111111101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7072|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfhax6_reg  (
    .a({open_n68601,_al_u7062_o}),
    .b({_al_u7071_o,_al_u6879_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [16],_al_u7072_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7072_o,open_n68619}),
    .q({open_n68623,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] }));  // ../RTL/cortexm0ds_logic.v(18495)
  // ../RTL/cortexm0ds_logic.v(18489)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*A*~(D*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(C*A*~(D*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0111111101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7075|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zdhax6_reg  (
    .a({open_n68624,_al_u7062_o}),
    .b({_al_u7074_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q7miu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [17],_al_u7075_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cmziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7075_o,open_n68642}),
    .q({open_n68646,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] }));  // ../RTL/cortexm0ds_logic.v(18489)
  // ../RTL/cortexm0ds_logic.v(18483)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*A*~(D*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(C*A*~(D*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0111111101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7078|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cchax6_reg  (
    .a({open_n68647,_al_u7062_o}),
    .b({_al_u7077_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R4miu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20],_al_u7078_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7078_o,open_n68665}),
    .q({open_n68669,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] }));  // ../RTL/cortexm0ds_logic.v(18483)
  // ../RTL/cortexm0ds_logic.v(18477)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*A*~(D*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("~(C*A*~(D*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111101011111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0111111101011111),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7081|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fahax6_reg  (
    .a({open_n68670,_al_u7062_o}),
    .b({_al_u7080_o,_al_u6926_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21],_al_u7081_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7081_o,open_n68688}),
    .q({open_n68692,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] }));  // ../RTL/cortexm0ds_logic.v(18477)
  // ../RTL/cortexm0ds_logic.v(18471)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~B*D)"),
    //.LUT1("(D*~(B*~(~C*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111111111),
    .INIT_LUT1(16'b0011011100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7083|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I8hax6_reg  (
    .a({_al_u6930_o,open_n68693}),
    .b({_al_u6941_o,_al_u7083_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vacow6 ,_al_u7085_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv ,_al_u7062_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7083_o,open_n68707}),
    .q({open_n68711,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] }));  // ../RTL/cortexm0ds_logic.v(18471)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~((D*B))*~(A)+C*(D*B)*~(A)+~(C)*(D*B)*A+C*(D*B)*A)"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0010011110101111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u7085|_al_u7084  (
    .a({open_n68712,_al_u4289_o}),
    .b({_al_u7084_o,_al_u4290_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [20]}),
    .f({_al_u7085_o,_al_u7084_o}));
  // ../RTL/cortexm0ds_logic.v(18085)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*A*~(D*~B))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111101011111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7088|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C37ax6_reg  (
    .a({open_n68733,_al_u7062_o}),
    .b({_al_u7087_o,_al_u6962_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24],_al_u7088_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7088_o,open_n68747}),
    .q({open_n68751,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] }));  // ../RTL/cortexm0ds_logic.v(18085)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7091|_al_u7090  (
    .b({open_n68754,_al_u604_o}),
    .c({_al_u7090_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hirpw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hvcow6_lutinv ,_al_u6842_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fucow6_lutinv ,_al_u7090_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(A)*~(C)+~(D*~B)*A*~(C)+~(~(D*~B))*A*C+~(D*~B)*A*C)"),
    //.LUT1("(D*C*~(B*~A))"),
    .INIT_LUT0(16'b1010110010101111),
    .INIT_LUT1(16'b1011000000000000),
    .MODE("LOGIC"))
    \_al_u7092|_al_u6839  (
    .a({_al_u6826_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh3ju6 }),
    .b({_al_u6836_o,_al_u6830_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fucow6_lutinv ,_al_u6838_o}),
    .f({_al_u7092_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxlow6_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~(~C*~B)*~(~D*~A))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~(~C*~B)*~(~D*~A))"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111110010101000),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111110010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7094|_al_u7093  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ,open_n68799}),
    .b({_al_u7093_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tucow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Piziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Alziu6 ,_al_u7090_o}),
    .f({_al_u7094_o,_al_u7093_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7096|_al_u7097  (
    .b({_al_u7094_o,_al_u7096_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjziu6 ,_al_u6930_o}),
    .f({_al_u7096_o,_al_u7097_o}));
  // ../RTL/cortexm0ds_logic.v(19759)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u709|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Do6bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[10] }),
    .mi({open_n68860,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,_al_u894_o}),
    .q({open_n68865,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[10] }));  // ../RTL/cortexm0ds_logic.v(19759)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*~B))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b0101000001000000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u7100|_al_u7101  (
    .a({open_n68866,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ,_al_u6846_o}),
    .c({_al_u6856_o,_al_u7100_o}),
    .d({_al_u7099_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }),
    .f({_al_u7100_o,_al_u7101_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*~(~C*A))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1111010111000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u7104|_al_u7103  (
    .a({open_n68887,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .b({_al_u7103_o,_al_u7093_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xv6ow6 }),
    .d({_al_u6870_o,_al_u6876_o}),
    .f({_al_u7104_o,_al_u7103_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~B)*~(~C*A))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~(~D*~B)*~(~C*A))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111010111000100),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111010111000100),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7108|_al_u7107  (
    .a({open_n68908,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .b({_al_u7093_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plcow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlcow6 }),
    .f({_al_u7108_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejcow6 }));
  // ../RTL/cortexm0ds_logic.v(17901)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*~D)"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("~(C*B*~D)"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100111111),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b1111111100111111),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u7109|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zazpw6_reg  (
    .b({_al_u7108_o,_al_u7109_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ,_al_u5911_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ukcow6 ,_al_u7092_o}),
    .f({_al_u7109_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .q({open_n68955,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[24] }));  // ../RTL/cortexm0ds_logic.v(17901)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~B)*~(~C*A))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~(~D*~B)*~(~C*A))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111010111000100),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b1111010111000100),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7112|_al_u7111  (
    .a({open_n68956,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .b({_al_u7093_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgcow6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iecow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahcow6 }),
    .f({_al_u7112_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iecow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*~B)*~(~D*~A))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1111110010101000),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u7116|_al_u7115  (
    .a({open_n68981,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3cow6 ,_al_u7093_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ,_al_u6952_o}),
    .d({_al_u6949_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G6cow6 }),
    .f({_al_u7116_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3cow6 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*~(~C*~A))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1111101011001000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u7120|_al_u7119  (
    .a({open_n69002,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0cow6 ,_al_u7093_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1cow6 }),
    .d({_al_u7119_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0cow6 }),
    .f({_al_u7120_o,_al_u7119_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~(D*~A)))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(C*~(D*~A)))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0100110000001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0100110000001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7122|_al_u7121  (
    .a({open_n69023,_al_u6913_o}),
    .b({open_n69024,_al_u7120_o}),
    .c({_al_u7121_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .d({_al_u7092_o,_al_u6925_o}),
    .f({_al_u7122_o,_al_u7121_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D*~A)))"),
    //.LUT1("(~(~D*~C)*~(~B*~A))"),
    .INIT_LUT0(16'b0100110000001100),
    .INIT_LUT1(16'b1110111011100000),
    .MODE("LOGIC"))
    \_al_u7124|_al_u7125  (
    .a({_al_u6822_o,_al_u6827_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kjziu6_lutinv ,_al_u7124_o}),
    .c({_al_u7093_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xbcow6_lutinv }),
    .d({_al_u6829_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iimow6 }),
    .f({_al_u7124_o,_al_u7125_o}));
  // ../RTL/cortexm0ds_logic.v(17905)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*~D)"),
    //.LUT1("(D*~(~C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100111111),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u7126|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yizpw6_reg  (
    .b({_al_u6820_o,_al_u7126_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlziu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbliu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u7125_o,_al_u7092_o}),
    .f({_al_u7126_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .q({open_n69087,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[29] }));  // ../RTL/cortexm0ds_logic.v(17905)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~D))"),
    //.LUT1("(D*~C*~B*A)"),
    .INIT_LUT0(16'b0000111100000011),
    .INIT_LUT1(16'b0000001000000000),
    .MODE("LOGIC"))
    \_al_u7129|_al_u7128  (
    .a({_al_u7128_o,open_n69088}),
    .b({_al_u3874_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uzaiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qaciu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzjpw6 ,_al_u3874_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ,_al_u7128_o}));
  // ../RTL/cortexm0ds_logic.v(17853)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u712|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsxpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M6kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxjpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[10] }),
    .mi({open_n69112,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ,_al_u892_o}),
    .q({open_n69128,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[10] }));  // ../RTL/cortexm0ds_logic.v(17853)
  // ../RTL/cortexm0ds_logic.v(18607)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(~(C*~B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0100010111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7130|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eliax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ,open_n69129}),
    .b({_al_u7128_o,_al_u7130_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] ,_al_u7131_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdspw6 ,_al_u7028_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7130_o,open_n69143}),
    .q({open_n69147,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[0] }));  // ../RTL/cortexm0ds_logic.v(18607)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7131|_al_u4295  (
    .b({open_n69150,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .c({_al_u4295_o,_al_u609_o}),
    .d({_al_u3874_o,_al_u1788_o}),
    .f({_al_u7131_o,_al_u4295_o}));
  // ../RTL/cortexm0ds_logic.v(18613)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(~(C*~B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0100010111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7133|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aniax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ,open_n69175}),
    .b({_al_u7128_o,_al_u7133_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] ,_al_u7131_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpmpw6 ,_al_u7032_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7133_o,open_n69189}),
    .q({open_n69193,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[2] }));  // ../RTL/cortexm0ds_logic.v(18613)
  // ../RTL/cortexm0ds_logic.v(17427)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(C*~B)*~(D*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(C*~B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0100010111001111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0100010111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7135|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qhmpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ,open_n69194}),
    .b({_al_u7128_o,_al_u7135_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] ,_al_u7131_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xiipw6 ,_al_u7036_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7135_o,open_n69212}),
    .q({open_n69216,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[3] }));  // ../RTL/cortexm0ds_logic.v(17427)
  // ../RTL/cortexm0ds_logic.v(18601)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(~(D*~B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0100110001011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7137|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ijiax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ,open_n69217}),
    .b({_al_u7128_o,_al_u7137_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2iax6 ,_al_u7131_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] ,_al_u7041_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7137_o,open_n69231}),
    .q({open_n69235,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[4] }));  // ../RTL/cortexm0ds_logic.v(18601)
  // ../RTL/cortexm0ds_logic.v(17295)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(D*~B)*~(C*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(D*~B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0100110001011111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0100110001011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7139|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbkpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ,open_n69236}),
    .b({_al_u7128_o,_al_u7139_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F4iax6 ,_al_u7131_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] ,_al_u7045_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7139_o,open_n69254}),
    .q({open_n69258,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[5] }));  // ../RTL/cortexm0ds_logic.v(17295)
  // ../RTL/cortexm0ds_logic.v(17605)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(C*~B)*~(D*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(C*~B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0100010111001111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0100010111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7141|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pcrpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xibiu6 ,open_n69259}),
    .b({_al_u7128_o,_al_u7141_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] ,_al_u7131_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5mpw6 ,_al_u7057_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7141_o,open_n69277}),
    .q({open_n69281,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_ipsr_o[1] }));  // ../RTL/cortexm0ds_logic.v(17605)
  // ../RTL/cortexm0ds_logic.v(19782)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7144|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq7bx6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u6985_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idkow6 ,_al_u7144_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7144_o,open_n69295}),
    .q({open_n69299,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] }));  // ../RTL/cortexm0ds_logic.v(19782)
  // ../RTL/cortexm0ds_logic.v(17238)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(~(~D*~A)*~(B)*~(C)+~(~D*~A)*B*~(C)+~(~(~D*~A))*B*C+~(~D*~A)*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b1100111111001010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7146|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bfjpw6_reg  (
    .a({_al_u6216_o,_al_u7092_o}),
    .b({_al_u2270_o,_al_u7117_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ,_al_u7146_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7146_o,open_n69312}),
    .q({open_n69316,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[2] }));  // ../RTL/cortexm0ds_logic.v(17238)
  // ../RTL/cortexm0ds_logic.v(17475)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b1111001111100010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7148|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Arnpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vioiu6_lutinv ,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ,_al_u7126_o}),
    .c({_al_u2281_o,_al_u7148_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5liu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7148_o,open_n69329}),
    .q({open_n69333,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[3] }));  // ../RTL/cortexm0ds_logic.v(17475)
  // ../RTL/cortexm0ds_logic.v(18555)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7151|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhax6_reg  (
    .a({_al_u7060_o,open_n69334}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7151_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0how6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3],_al_u7032_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7151_o,open_n69352}),
    .q({open_n69356,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] }));  // ../RTL/cortexm0ds_logic.v(18555)
  // ../RTL/cortexm0ds_logic.v(18549)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7154|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwhax6_reg  (
    .a({_al_u7060_o,open_n69357}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7154_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rwgow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4],_al_u7036_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7154_o,open_n69375}),
    .q({open_n69379,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] }));  // ../RTL/cortexm0ds_logic.v(18549)
  // ../RTL/cortexm0ds_logic.v(18543)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7157|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vuhax6_reg  (
    .a({_al_u7060_o,open_n69380}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7157_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkfow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5],_al_u7041_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7157_o,open_n69398}),
    .q({open_n69402,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] }));  // ../RTL/cortexm0ds_logic.v(18543)
  // ../RTL/cortexm0ds_logic.v(18825)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u715|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5qax6_reg  (
    .a({_al_u705_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv9pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u711_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u714_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[0] }),
    .mi({open_n69406,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yv9pw6 }),
    .q({open_n69422,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[0] }));  // ../RTL/cortexm0ds_logic.v(18825)
  // ../RTL/cortexm0ds_logic.v(18537)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7160|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zshax6_reg  (
    .a({_al_u7060_o,open_n69423}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7160_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xneow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6],_al_u7045_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7160_o,open_n69437}),
    .q({open_n69441,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] }));  // ../RTL/cortexm0ds_logic.v(18537)
  // ../RTL/cortexm0ds_logic.v(17611)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7163|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lerpw6_reg  (
    .a({_al_u7060_o,open_n69442}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7163_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr6ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2],_al_u7057_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7163_o,open_n69456}),
    .q({open_n69460,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }));  // ../RTL/cortexm0ds_logic.v(17611)
  // ../RTL/cortexm0ds_logic.v(17961)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7166|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A32qw6_reg  (
    .a({_al_u7060_o,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7117_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M2cow6 ,_al_u7166_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7166_o,open_n69474}),
    .q({open_n69478,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] }));  // ../RTL/cortexm0ds_logic.v(17961)
  // ../RTL/cortexm0ds_logic.v(17955)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7169|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D12qw6_reg  (
    .a({_al_u7060_o,open_n69479}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7169_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qxbow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29],_al_u7122_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7169_o,open_n69493}),
    .q({open_n69497,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] }));  // ../RTL/cortexm0ds_logic.v(17955)
  // ../RTL/cortexm0ds_logic.v(17729)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7172|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Awupw6_reg  (
    .a({_al_u7060_o,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7126_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ow6 ,_al_u7172_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7172_o,open_n69515}),
    .q({open_n69519,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] }));  // ../RTL/cortexm0ds_logic.v(17729)
  // ../RTL/cortexm0ds_logic.v(19926)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7175|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P7bbx6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u6981_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A0mow6 ,_al_u7175_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7175_o,open_n69537}),
    .q({open_n69541,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] }));  // ../RTL/cortexm0ds_logic.v(19926)
  // ../RTL/cortexm0ds_logic.v(19741)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7178|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J06bx6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u6989_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdjow6 ,_al_u7178_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7178_o,open_n69559}),
    .q({open_n69563,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] }));  // ../RTL/cortexm0ds_logic.v(19741)
  // ../RTL/cortexm0ds_logic.v(19734)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7181|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mw5bx6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u6994_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eriow6 ,_al_u7181_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7181_o,open_n69581}),
    .q({open_n69585,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] }));  // ../RTL/cortexm0ds_logic.v(19734)
  // ../RTL/cortexm0ds_logic.v(18525)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7184|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hphax6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u6998_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvdow6 ,_al_u7184_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7184_o,open_n69599}),
    .q({open_n69603,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] }));  // ../RTL/cortexm0ds_logic.v(18525)
  // ../RTL/cortexm0ds_logic.v(18519)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7187|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Knhax6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7002_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Prdow6 ,_al_u7187_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7187_o,open_n69621}),
    .q({open_n69625,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] }));  // ../RTL/cortexm0ds_logic.v(18519)
  // ../RTL/cortexm0ds_logic.v(18513)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7190|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlhax6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7006_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hndow6 ,_al_u7190_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7190_o,open_n69639}),
    .q({open_n69643,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] }));  // ../RTL/cortexm0ds_logic.v(18513)
  // ../RTL/cortexm0ds_logic.v(18507)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7193|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjhax6_reg  (
    .a({_al_u7060_o,_al_u6969_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7010_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eidow6 ,_al_u7193_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7193_o,open_n69661}),
    .q({open_n69665,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] }));  // ../RTL/cortexm0ds_logic.v(18507)
  // ../RTL/cortexm0ds_logic.v(17245)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b1111001111100010),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b1111001111100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7195|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qijpw6_reg  (
    .a({_al_u6236_o,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ,_al_u7097_o}),
    .c({_al_u2429_o,_al_u7195_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7195_o,open_n69682}),
    .q({open_n69686,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[1] }));  // ../RTL/cortexm0ds_logic.v(17245)
  // ../RTL/cortexm0ds_logic.v(18531)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7198|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drhax6_reg  (
    .a({_al_u7060_o,open_n69687}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7198_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dkeow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7],_al_u7049_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7198_o,open_n69701}),
    .q({open_n69705,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] }));  // ../RTL/cortexm0ds_logic.v(18531)
  // ../RTL/cortexm0ds_logic.v(17716)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7201|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Equpw6_reg  (
    .a({_al_u7060_o,open_n69706}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7201_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W48ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8],_al_u7053_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7201_o,open_n69720}),
    .q({open_n69724,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] }));  // ../RTL/cortexm0ds_logic.v(17716)
  // ../RTL/cortexm0ds_logic.v(17259)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7204|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqjpw6_reg  (
    .a({_al_u7060_o,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7097_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfziu6 ,_al_u7204_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7204_o,open_n69738}),
    .q({open_n69742,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] }));  // ../RTL/cortexm0ds_logic.v(17259)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~(D*C)*~(~B*A))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~(D*C)*~(~B*A))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000110111011101),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7206|_al_u2797  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 ,open_n69743}),
    .b({_al_u1299_o,_al_u1299_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Et8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ubypw6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjoiu6 }),
    .f({_al_u7206_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(17322)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D*~A)))"),
    //.LUT1("(C*~(~D*~(B*~A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000011100000011),
    .INIT_LUT1(16'b1111000001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7207|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pzkpw6_reg  (
    .a({_al_u7013_o,_al_u7101_o}),
    .b({_al_u7027_o,_al_u7207_o}),
    .c({_al_u7206_o,_al_u7208_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nn8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u4172_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7207_o,open_n69780}),
    .q({open_n69784,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_tbit_o }));  // ../RTL/cortexm0ds_logic.v(17322)
  // ../RTL/cortexm0ds_logic.v(18465)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7211|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6hax6_reg  (
    .a({_al_u7060_o,open_n69785}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7211_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lqcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25],_al_u7101_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7211_o,open_n69803}),
    .q({open_n69807,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] }));  // ../RTL/cortexm0ds_logic.v(18465)
  // ../RTL/cortexm0ds_logic.v(18459)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7214|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4hax6_reg  (
    .a({_al_u7060_o,open_n69808}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7214_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rmcow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26],_al_u7105_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7214_o,open_n69826}),
    .q({open_n69830,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] }));  // ../RTL/cortexm0ds_logic.v(18459)
  // ../RTL/cortexm0ds_logic.v(18453)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~(B*~A)))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011111100001111),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7217|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R2hax6_reg  (
    .a({_al_u7060_o,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7109_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vhcow6 ,_al_u7217_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7217_o,open_n69844}),
    .q({open_n69848,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] }));  // ../RTL/cortexm0ds_logic.v(18453)
  // ../RTL/cortexm0ds_logic.v(18816)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u721|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Enpax6_reg  (
    .a({_al_u717_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u718_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u719_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u720_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] }),
    .mi({open_n69852,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ib0iu6 ,_al_u717_o}),
    .q({open_n69868,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] }));  // ../RTL/cortexm0ds_logic.v(18816)
  // ../RTL/cortexm0ds_logic.v(18447)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~(B*~A)))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("~(C*~(D*~(B*~A)))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111100001111),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b1011111100001111),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7220|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0hax6_reg  (
    .a({_al_u7060_o,_al_u7092_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Egziu6 ,_al_u7113_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zccow6 ,_al_u7220_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgziu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7220_o,open_n69886}),
    .q({open_n69890,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] }));  // ../RTL/cortexm0ds_logic.v(18447)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*D))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(~C*~(B*D))"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b0000001100001111),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0000001100001111),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7223|_al_u7222  (
    .b({_al_u2420_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P9niu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .d({_al_u7222_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv }),
    .f({_al_u7223_o,_al_u7222_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u7224|_al_u2799  (
    .b({_al_u6242_o,open_n69919}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv }),
    .d({_al_u7223_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ph8iu6_lutinv }),
    .f({_al_u7224_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ug8iu6_lutinv }));
  // ../RTL/cortexm0ds_logic.v(20165)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~A)))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~(B*~(D*~A)))"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000011100000011),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u7225|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5ibx6_reg  (
    .a({open_n69940,_al_u7122_o}),
    .b({open_n69941,_al_u7224_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] ,_al_u7225_o}),
    .clk(XTAL1_wire),
    .d({_al_u7222_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yi8iu6_lutinv }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u7225_o,open_n69959}),
    .q({open_n69963,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_apsr_o[0] }));  // ../RTL/cortexm0ds_logic.v(20165)
  // ../RTL/cortexm0ds_logic.v(18815)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u727|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elpax6_reg  (
    .a({_al_u723_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A59pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u725_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u726_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[13] }),
    .mi({open_n69974,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bb0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A59pw6 }),
    .q({open_n69979,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] }));  // ../RTL/cortexm0ds_logic.v(18815)
  // ../RTL/cortexm0ds_logic.v(18814)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u733|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejpax6_reg  (
    .a({_al_u729_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv8pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u731_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u732_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] }),
    .mi({open_n69990,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ua0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wv8pw6 }),
    .q({open_n69995,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[14] }));  // ../RTL/cortexm0ds_logic.v(18814)
  // ../RTL/cortexm0ds_logic.v(19794)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u739|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zb8bx6_reg  (
    .a({_al_u735_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u736_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u737_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u738_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[15] }),
    .mi({open_n69999,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Na0iu6 ,_al_u735_o}),
    .q({open_n70015,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[15] }));  // ../RTL/cortexm0ds_logic.v(19794)
  // ../RTL/cortexm0ds_logic.v(18812)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u751|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Efpax6_reg  (
    .a({_al_u747_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W38pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u749_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u750_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[17] }),
    .mi({open_n70019,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z90iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W38pw6 }),
    .q({open_n70035,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] }));  // ../RTL/cortexm0ds_logic.v(18812)
  // ../RTL/cortexm0ds_logic.v(18811)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u757|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Edpax6_reg  (
    .a({_al_u753_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u754_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u755_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u756_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] }),
    .mi({open_n70046,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S90iu6 ,_al_u753_o}),
    .q({open_n70051,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[18] }));  // ../RTL/cortexm0ds_logic.v(18811)
  // ../RTL/cortexm0ds_logic.v(18810)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u763|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ebpax6_reg  (
    .a({_al_u759_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u760_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u761_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u762_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] }),
    .mi({open_n70062,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L90iu6 ,_al_u760_o}),
    .q({open_n70067,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] }));  // ../RTL/cortexm0ds_logic.v(18810)
  // ../RTL/cortexm0ds_logic.v(19722)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u769|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq5bx6_reg  (
    .a({_al_u765_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({_al_u766_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({_al_u767_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u768_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] }),
    .mi({open_n70078,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E90iu6 ,_al_u767_o}),
    .q({open_n70083,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[1] }));  // ../RTL/cortexm0ds_logic.v(19722)
  // ../RTL/cortexm0ds_logic.v(17451)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u775|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E7npw6_reg  (
    .a({_al_u771_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({_al_u772_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L27pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u774_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] }),
    .mi({open_n70094,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X80iu6 ,_al_u772_o}),
    .q({open_n70099,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] }));  // ../RTL/cortexm0ds_logic.v(17451)
  // ../RTL/cortexm0ds_logic.v(17450)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u781|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5npw6_reg  (
    .a({_al_u777_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({_al_u778_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({_al_u779_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u780_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] }),
    .mi({open_n70110,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q80iu6 ,_al_u780_o}),
    .q({open_n70115,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[21] }));  // ../RTL/cortexm0ds_logic.v(17450)
  // ../RTL/cortexm0ds_logic.v(20007)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u787|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T7fbx6_reg  (
    .a({_al_u783_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ml6pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u786_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[22] }),
    .mi({open_n70126,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J80iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6pw6 }),
    .q({open_n70131,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] }));  // ../RTL/cortexm0ds_logic.v(20007)
  // ../RTL/cortexm0ds_logic.v(18066)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u793|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gt6ax6_reg  (
    .a({_al_u789_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({_al_u790_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Za6pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u792_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] }),
    .mi({open_n70142,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C80iu6 ,_al_u790_o}),
    .q({open_n70147,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[23] }));  // ../RTL/cortexm0ds_logic.v(18066)
  // ../RTL/cortexm0ds_logic.v(18802)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u799|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fvoax6_reg  (
    .a({_al_u795_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u796_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u797_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u798_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] }),
    .mi({open_n70151,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V70iu6 ,_al_u795_o}),
    .q({open_n70167,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] }));  // ../RTL/cortexm0ds_logic.v(18802)
  // ../RTL/cortexm0ds_logic.v(18807)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u805|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E5pax6_reg  (
    .a({_al_u801_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({_al_u802_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs5pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u804_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[25] }),
    .mi({open_n70178,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O70iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs5pw6 }),
    .q({open_n70183,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[25] }));  // ../RTL/cortexm0ds_logic.v(18807)
  // ../RTL/cortexm0ds_logic.v(18831)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u811|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vgqax6_reg  (
    .a({_al_u807_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({_al_u808_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({_al_u809_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wk5pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] }),
    .mi({open_n70194,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H70iu6 ,_al_u809_o}),
    .q({open_n70199,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[26] }));  // ../RTL/cortexm0ds_logic.v(18831)
  // ../RTL/cortexm0ds_logic.v(18804)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u817|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzoax6_reg  (
    .a({_al_u813_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u814_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u815_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u816_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] }),
    .mi({open_n70210,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A70iu6 ,_al_u813_o}),
    .q({open_n70215,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[27] }));  // ../RTL/cortexm0ds_logic.v(18804)
  // ../RTL/cortexm0ds_logic.v(20167)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u823|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7ibx6_reg  (
    .a({_al_u819_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F15pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u821_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u822_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[28] }),
    .mi({open_n70219,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({_al_u823_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F15pw6 }),
    .q({open_n70235,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[28] }));  // ../RTL/cortexm0ds_logic.v(20167)
  // ../RTL/cortexm0ds_logic.v(17538)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u829|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhppw6_reg  (
    .a({_al_u825_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rt4pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u828_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[29] }),
    .mi({open_n70246,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M60iu6 ,_al_u825_o}),
    .q({open_n70251,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[29] }));  // ../RTL/cortexm0ds_logic.v(17538)
  // ../RTL/cortexm0ds_logic.v(18795)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u835|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khoax6_reg  (
    .a({_al_u831_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u832_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({_al_u833_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[30] }),
    .mi({open_n70262,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50iu6 ,_al_u832_o}),
    .q({open_n70267,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] }));  // ../RTL/cortexm0ds_logic.v(18795)
  // ../RTL/cortexm0ds_logic.v(17642)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u841|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7spw6_reg  (
    .a({_al_u837_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ha4pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({_al_u839_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u840_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] }),
    .mi({open_n70271,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P40iu6 ,_al_u837_o}),
    .q({open_n70287,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[6] }));  // ../RTL/cortexm0ds_logic.v(17642)
  // ../RTL/cortexm0ds_logic.v(17945)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u847|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jp1qw6_reg  (
    .a({_al_u843_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({_al_u844_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D14pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u846_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] }),
    .mi({open_n70298,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U30iu6 ,_al_u844_o}),
    .q({open_n70303,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[9] }));  // ../RTL/cortexm0ds_logic.v(17945)
  // ../RTL/cortexm0ds_logic.v(18824)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u853|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A3qax6_reg  (
    .a({_al_u849_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({_al_u850_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({_al_u851_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u852_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] }),
    .mi({open_n70314,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R50iu6 ,_al_u851_o}),
    .q({open_n70319,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] }));  // ../RTL/cortexm0ds_logic.v(18824)
  // ../RTL/cortexm0ds_logic.v(17543)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u859|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lrppw6_reg  (
    .a({_al_u855_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5pow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A4pow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u858_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] }),
    .mi({open_n70323,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D50iu6 ,_al_u855_o}),
    .q({open_n70339,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] }));  // ../RTL/cortexm0ds_logic.v(17543)
  // ../RTL/cortexm0ds_logic.v(18923)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u865|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjvax6_reg  (
    .a({_al_u861_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({_al_u862_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0pow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u864_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] }),
    .mi({open_n70350,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F60iu6 ,_al_u862_o}),
    .q({open_n70355,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[2] }));  // ../RTL/cortexm0ds_logic.v(18923)
  // ../RTL/cortexm0ds_logic.v(17535)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u871|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbppw6_reg  (
    .a({_al_u867_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({_al_u868_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({_al_u869_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u870_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] }),
    .mi({open_n70366,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K50iu6 ,_al_u867_o}),
    .q({open_n70371,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[3] }));  // ../RTL/cortexm0ds_logic.v(17535)
  // ../RTL/cortexm0ds_logic.v(18976)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u877|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S7yax6_reg  (
    .a({_al_u873_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({_al_u874_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({_al_u875_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u876_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[5] }),
    .mi({open_n70382,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W40iu6 ,_al_u875_o}),
    .q({open_n70387,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[5] }));  // ../RTL/cortexm0ds_logic.v(18976)
  // ../RTL/cortexm0ds_logic.v(18819)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u883|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dtpax6_reg  (
    .a({_al_u879_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({_al_u880_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhoow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u882_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[8] }),
    .mi({open_n70398,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B40iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhoow6 }),
    .q({open_n70403,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[8] }));  // ../RTL/cortexm0ds_logic.v(18819)
  // ../RTL/cortexm0ds_logic.v(19717)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u889|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Og5bx6_reg  (
    .a({_al_u885_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({_al_u886_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({_al_u887_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u888_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[7] }),
    .mi({open_n70407,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I40iu6 ,_al_u887_o}),
    .q({open_n70423,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[7] }));  // ../RTL/cortexm0ds_logic.v(19717)
  // ../RTL/cortexm0ds_logic.v(18920)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u895|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vdvax6_reg  (
    .a({_al_u891_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({_al_u892_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cenow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u894_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] }),
    .mi({open_n70427,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wb0iu6 ,_al_u891_o}),
    .q({open_n70443,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[10] }));  // ../RTL/cortexm0ds_logic.v(18920)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u901|_al_u902  (
    .a({_al_u897_o,open_n70444}),
    .b({_al_u898_o,open_n70445}),
    .c({_al_u899_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 }),
    .d({_al_u900_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xuzhu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pb0iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [11]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u907|_al_u904  (
    .c({_al_u906_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxupw6 }),
    .d({_al_u904_o,_al_u903_o}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ,_al_u904_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(D*C))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~B*~A*~(D*C))"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000100010001),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000100010001),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u910|_al_u4164  (
    .a({open_n70498,_al_u908_o}),
    .b({_al_u908_o,_al_u3591_o}),
    .c({_al_u909_o,_al_u607_o}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F85iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vo3ju6_lutinv }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 ,_al_u4164_o}));
  // ../RTL/cortexm0ds_logic.v(17444)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*~B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(D*C*~B*A)"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111111111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1101111111111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u913|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6_reg  (
    .a({open_n70523,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpyiu6 }),
    .b({open_n70524,_al_u913_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0kax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aj1ju6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O25iu6 ),
    .clk(XTAL1_wire),
    .d({_al_u912_o,_al_u920_o}),
    .f({_al_u913_o,open_n70542}),
    .q({open_n70546,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Htmpw6 }));  // ../RTL/cortexm0ds_logic.v(17444)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u920|_al_u2749  (
    .a({_al_u696_o,_al_u696_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A95iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Irmpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iekax6 }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oikax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfspw6 }),
    .f({_al_u920_o,_al_u2749_o}));
  // ../RTL/cortexm0ds_logic.v(18405)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u923|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 ,open_n70573}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u923_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 }),
    .q({open_n70590,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydgax6 }));  // ../RTL/cortexm0ds_logic.v(18405)
  // ../RTL/cortexm0ds_logic.v(18250)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u924|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ,open_n70591}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 ,open_n70592}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H0ebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u924_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 }),
    .q({open_n70609,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 }));  // ../RTL/cortexm0ds_logic.v(18250)
  // ../RTL/cortexm0ds_logic.v(18043)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u925|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6_reg  (
    .a({_al_u923_o,open_n70610}),
    .b({_al_u924_o,open_n70611}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .f({_al_u925_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .q({open_n70632,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym3qw6 }));  // ../RTL/cortexm0ds_logic.v(18043)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u933|_al_u931  (
    .b({_al_u932_o,_al_u930_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T1vpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufopw6 }),
    .d({_al_u931_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qyniu6_lutinv }),
    .f({_al_u933_o,_al_u931_o}));
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~(C*B)))"),
    //.LUT1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000010101010),
    .INIT_LUT1(16'b1010100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u935|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b7  (
    .a({_al_u470_o,_al_u3370_o}),
    .b({b_pad_gpio_porta_pad[7],\u_cmsdk_mcu/HWDATA [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qo3bx6 }),
    .mi({open_n70665,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u935_o,_al_u3371_o}),
    .q({open_n70669,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]}));  // ../RTL/gpio_apbif.v(262)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(B*A)))"),
    //.LUTF1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("(~C*~(D*~(B*A)))"),
    //.LUTG1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001111),
    .INIT_LUTF1(16'b1100100000001000),
    .INIT_LUTG0(16'b0000100000001111),
    .INIT_LUTG1(16'b1100100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u937|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [7],\u_cmsdk_mcu/HWDATA [7]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [7],_al_u3072_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [7]}),
    .mi({open_n70673,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [7],_al_u3073_o}),
    .q({open_n70688,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7]}));  // ../RTL/gpio_apbif.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~B*C*~D+~A*~B*C*D+~A*B*C*D)"),
    //.LUTF1("(~D*~C*~(~B*A))"),
    //.LUTG0("(~A*~B*C*~D+~A*~B*C*D+~A*B*C*D)"),
    //.LUTG1("(~D*~C*~(~B*A))"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000000001101),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000000001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u938|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b2_rom0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .f({_al_u938_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [2]}));
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D*~C*~A))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(D*~C*~A))"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011011100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0011011100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u939|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b7  (
    .a({open_n70713,_al_u939_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [7],_al_u946_o}),
    .c({_al_u938_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u935_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u939_o,open_n70730}),
    .q({open_n70734,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [7]}));  // ../RTL/gpio_apbif.v(453)
  EG_PHY_PAD #(
    //.LOCATION("T4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u94 (
    .ipad(NRST),
    .di(NRST_pad));  // ../RTL/M0demo.v(7)
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011111111110101),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011111111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u940|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [7],open_n70752}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [7],open_n70753}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2494_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n70757,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u940_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n113 }),
    .q({open_n70772,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [7]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_apbif.v(343)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u941|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [7],open_n70773}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [7],open_n70774}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2496_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n70785,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u941_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n68 }),
    .q({open_n70789,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [7]}));  // ../RTL/gpio_apbif.v(343)
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C@D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(C@D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u942|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b7  (
    .c({_al_u941_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [7]}),
    .clk(1'b1),
    .d({_al_u940_o,b_pad_gpio_porta_pad[7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u942_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [7]}),
    .q({open_n70814,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [7]}));  // ../RTL/gpio_ctrl.v(184)
  // ../RTL/gpio_apbif.v(242)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000010101100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u943|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7],open_n70815}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7],open_n70816}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2490_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n70827,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b7/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n203 }),
    .q({open_n70831,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [7]}));  // ../RTL/gpio_apbif.v(242)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b1010111111110011),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1010111111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u944|_al_u945  (
    .a({_al_u942_o,open_n70832}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b7/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,_al_u467_o}),
    .f({_al_u944_o,_al_u945_o}));
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~A*~((C*B))*~(D)+~A*(C*B)*~(D)+~(~A)*(C*B)*D+~A*(C*B)*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~A*~((C*B))*~(D)+~A*(C*B)*~(D)+~(~A)*(C*B)*D+~A*(C*B)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011111110101010),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u946|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b7  (
    .a({_al_u944_o,open_n70857}),
    .b({_al_u945_o,open_n70858}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [7],_al_u2492_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({open_n70862,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u946_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n158 }),
    .q({open_n70877,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [7]}));  // ../RTL/gpio_apbif.v(383)
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~(C*B)))"),
    //.LUTF1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTG0("(A*~(D*~(C*B)))"),
    //.LUTG1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000010101010),
    .INIT_LUTF1(16'b1010100000001000),
    .INIT_LUTG0(16'b1000000010101010),
    .INIT_LUTG1(16'b1010100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u948|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b6  (
    .a({_al_u470_o,_al_u3360_o}),
    .b({b_pad_gpio_porta_pad[6],\u_cmsdk_mcu/HWDATA [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lr9bx6 }),
    .mi({open_n70881,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u948_o,_al_u3361_o}),
    .q({open_n70896,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]}));  // ../RTL/gpio_apbif.v(262)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u95 (
    .do({open_n70898,open_n70899,open_n70900,\u_cmsdk_mcu/p0_out [15]}),
    .ts(\u_cmsdk_mcu/p0_outen [15]),
    .opad(P0[15]));  // ../RTL/cmsdk_mcu_pin_mux.v(141)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(B*A)))"),
    //.LUTF1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("(~C*~(D*~(B*A)))"),
    //.LUTG1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001111),
    .INIT_LUTF1(16'b1100100000001000),
    .INIT_LUTG0(16'b0000100000001111),
    .INIT_LUTG1(16'b1100100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u950|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [6],\u_cmsdk_mcu/HWDATA [6]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [6],_al_u3067_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [6]}),
    .mi({open_n70916,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [6],_al_u3068_o}),
    .q({open_n70931,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6]}));  // ../RTL/gpio_apbif.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~(~B*A))"),
    //.LUTF1("(~D*~C*~(~B*A))"),
    //.LUTG0("(~D*~C*~(~B*A))"),
    //.LUTG1("(~D*~C*~(~B*A))"),
    .INIT_LUTF0(16'b0000000000001101),
    .INIT_LUTF1(16'b0000000000001101),
    .INIT_LUTG0(16'b0000000000001101),
    .INIT_LUTG1(16'b0000000000001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u951|_al_u999  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .f({_al_u951_o,_al_u999_o}));
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    //.LUT1("(~D*~(~A*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000001111),
    .INIT_LUT1(16'b0000000011101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u952|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b6  (
    .a({_al_u948_o,open_n70956}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [6],open_n70957}),
    .c({_al_u951_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [6]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,b_pad_gpio_porta_pad[6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u952_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [6]}),
    .q({open_n70974,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [6]}));  // ../RTL/gpio_ctrl.v(184)
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~A*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u953|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b6  (
    .a({_al_u952_o,open_n70975}),
    .b({_al_u945_o,open_n70976}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [6],_al_u2492_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n70987,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u953_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n156 }),
    .q({open_n70991,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [6]}));  // ../RTL/gpio_apbif.v(383)
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u954|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [6],open_n70992}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [6],open_n70993}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2494_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n71004,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u954_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n111 }),
    .q({open_n71008,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [6]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_apbif.v(343)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u955|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [6],open_n71009}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [6],open_n71010}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2496_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n71021,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u955_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n66 }),
    .q({open_n71025,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [6]}));  // ../RTL/gpio_apbif.v(343)
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u956|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b6  (
    .b({_al_u954_o,_al_u956_o}),
    .c({_al_u955_o,_al_u958_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u566_o,_al_u953_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u956_o,open_n71040}),
    .q({open_n71044,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [6]}));  // ../RTL/gpio_apbif.v(453)
  // ../RTL/gpio_apbif.v(242)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000010101100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u957|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b6  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6],open_n71045}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6],open_n71046}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2490_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({open_n71057,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b6/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n201 }),
    .q({open_n71061,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [6]}));  // ../RTL/gpio_apbif.v(242)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u96 (
    .do({open_n71063,open_n71064,open_n71065,\u_cmsdk_mcu/p0_out [14]}),
    .ts(\u_cmsdk_mcu/p0_outen [14]),
    .opad(P0[14]));  // ../RTL/cmsdk_mcu_pin_mux.v(140)
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTF1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUTG1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000001110111),
    .INIT_LUTF1(16'b1010100000001000),
    .INIT_LUTG0(16'b0010000001110111),
    .INIT_LUTG1(16'b1010100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u960|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b5  (
    .a({_al_u470_o,\u_cmsdk_mcu/HWDATA [5]}),
    .b({b_pad_gpio_porta_pad[5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mk3bx6 }),
    .mi({open_n71081,\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u960_o,_al_u3279_o}),
    .q({open_n71096,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]}));  // ../RTL/gpio_apbif.v(262)
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b1100100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u962|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [5],\u_cmsdk_mcu/HWDATA [5]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [5],_al_u3062_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [5]}),
    .mi({open_n71107,\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [5],_al_u3063_o}),
    .q({open_n71111,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5]}));  // ../RTL/gpio_apbif.v(303)
  // ../RTL/gpio_apbif.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*~C*~(~B*A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*~C*~(~B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001101),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u963|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg3_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5],open_n71112}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,open_n71113}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,_al_u2496_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n52 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/HWDATA [5]}),
    .mi({open_n71117,\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u963_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n64 }),
    .q({open_n71132,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5]}));  // ../RTL/gpio_apbif.v(323)
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~D*~(~A*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u964|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b5  (
    .a({_al_u960_o,open_n71133}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [5],open_n71134}),
    .c({_al_u963_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,_al_u3063_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u964_o,open_n71148}),
    .q({open_n71152,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [5]}));  // ../RTL/gpio_ctrl.v(248)
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~A*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u965|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b5  (
    .a({_al_u964_o,open_n71153}),
    .b({_al_u945_o,open_n71154}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [5],_al_u2490_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/HWDATA [5]}),
    .mi({open_n71165,\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u965_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n199 }),
    .q({open_n71169,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [5]}));  // ../RTL/gpio_apbif.v(383)
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u966|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [5],open_n71170}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [5],open_n71171}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2492_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [5]}),
    .mi({open_n71182,\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u966_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n154 }),
    .q({open_n71186,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [5]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_apbif.v(343)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111001101011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u967|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [5],open_n71187}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [5],open_n71188}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2494_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [5]}),
    .mi({open_n71192,\u_cmsdk_mcu/HWDATA [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u967_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n109 }),
    .q({open_n71207,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [5]}));  // ../RTL/gpio_apbif.v(343)
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u968|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b5  (
    .b({_al_u966_o,_al_u968_o}),
    .c({_al_u967_o,_al_u970_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u566_o,_al_u965_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u968_o,open_n71222}),
    .q({open_n71226,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [5]}));  // ../RTL/gpio_apbif.v(453)
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    //.LUT1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000001111),
    .INIT_LUT1(16'b0000000010101100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u969|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5],open_n71227}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5],open_n71228}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [5]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,b_pad_gpio_porta_pad[5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b5/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [5]}),
    .q({open_n71245,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [5]}));  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u97 (
    .do({open_n71247,open_n71248,open_n71249,\u_cmsdk_mcu/p0_out [13]}),
    .ts(\u_cmsdk_mcu/p0_outen [13]),
    .opad(P0[13]));  // ../RTL/cmsdk_mcu_pin_mux.v(139)
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUT1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000001110111),
    .INIT_LUT1(16'b1010100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u972|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b4  (
    .a({_al_u470_o,\u_cmsdk_mcu/HWDATA [4]}),
    .b({b_pad_gpio_porta_pad[4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gihbx6 }),
    .mi({open_n71272,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u972_o,_al_u3274_o}),
    .q({open_n71276,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]}));  // ../RTL/gpio_apbif.v(262)
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b1100100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u974|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [4],\u_cmsdk_mcu/HWDATA [4]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [4],_al_u3057_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [4]}),
    .mi({open_n71287,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [4],_al_u3058_o}),
    .q({open_n71291,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4]}));  // ../RTL/gpio_apbif.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~(~B*A))"),
    //.LUT1("(~D*~C*~(~B*A))"),
    .INIT_LUT0(16'b0000000000001101),
    .INIT_LUT1(16'b0000000000001101),
    .MODE("LOGIC"))
    \_al_u975|_al_u987  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4:3]),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .f({_al_u975_o,_al_u987_o}));
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C@D)"),
    //.LUTF1("(~D*~(~A*~(C*B)))"),
    //.LUTG0("~(C@D)"),
    //.LUTG1("(~D*~(~A*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000001111),
    .INIT_LUTF1(16'b0000000011101010),
    .INIT_LUTG0(16'b1111000000001111),
    .INIT_LUTG1(16'b0000000011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u976|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b4  (
    .a({_al_u972_o,open_n71312}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [4],open_n71313}),
    .c({_al_u975_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [4]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,b_pad_gpio_porta_pad[4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u976_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [4]}),
    .q({open_n71334,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [4]}));  // ../RTL/gpio_ctrl.v(184)
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~A*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u977|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b4  (
    .a({_al_u976_o,open_n71335}),
    .b({_al_u945_o,open_n71336}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [4],_al_u2490_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/HWDATA [4]}),
    .mi({open_n71347,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u977_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n197 }),
    .q({open_n71351,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [4]}));  // ../RTL/gpio_apbif.v(383)
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011111111110101),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011111111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u978|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [4],open_n71352}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [4],open_n71353}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2492_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [4]}),
    .mi({open_n71357,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u978_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n152 }),
    .q({open_n71372,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [4]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_apbif.v(343)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u979|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [4],open_n71373}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [4],open_n71374}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2494_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [4]}),
    .mi({open_n71385,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u979_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n107 }),
    .q({open_n71389,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [4]}));  // ../RTL/gpio_apbif.v(343)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u98 (
    .do({open_n71391,open_n71392,open_n71393,\u_cmsdk_mcu/p0_out [12]}),
    .ts(\u_cmsdk_mcu/p0_outen [12]),
    .opad(P0[12]));  // ../RTL/cmsdk_mcu_pin_mux.v(138)
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u980|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b4  (
    .b({_al_u978_o,_al_u980_o}),
    .c({_al_u979_o,_al_u982_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u566_o,_al_u977_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u980_o,open_n71424}),
    .q({open_n71428,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [4]}));  // ../RTL/gpio_apbif.v(453)
  // ../RTL/gpio_apbif.v(242)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000010101100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u981|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4],open_n71429}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4],open_n71430}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2488_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [4]}),
    .mi({open_n71441,\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b4/B1_0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n242 }),
    .q({open_n71445,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [4]}));  // ../RTL/gpio_apbif.v(242)
  // ../RTL/gpio_apbif.v(262)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*C*D)"),
    //.LUT1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000001110111),
    .INIT_LUT1(16'b1010100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u984|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg0_b3  (
    .a({_al_u470_o,\u_cmsdk_mcu/HWDATA [3]}),
    .b({b_pad_gpio_porta_pad[3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n43 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Muhbx6 }),
    .mi({open_n71456,\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u984_o,_al_u3268_o}),
    .q({open_n71460,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]}));  // ../RTL/gpio_apbif.v(262)
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(B*A)))"),
    //.LUTF1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("(~C*~(D*~(B*A)))"),
    //.LUTG1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001111),
    .INIT_LUTF1(16'b1100100000001000),
    .INIT_LUTG0(16'b0000100000001111),
    .INIT_LUTG1(16'b1100100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u986|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [3],\u_cmsdk_mcu/HWDATA [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [3],_al_u3052_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [3]}),
    .mi({open_n71464,\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [3],_al_u3053_o}),
    .q({open_n71479,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3]}));  // ../RTL/gpio_apbif.v(303)
  // ../RTL/gpio_ctrl.v(184)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C@D)"),
    //.LUTF1("(~D*~(~A*~(C*B)))"),
    //.LUTG0("~(C@D)"),
    //.LUTG1("(~D*~(~A*~(C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000001111),
    .INIT_LUTF1(16'b0000000011101010),
    .INIT_LUTG0(16'b1111000000001111),
    .INIT_LUTG1(16'b0000000011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u988|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg0_b3  (
    .a({_al_u984_o,open_n71480}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [3],open_n71481}),
    .c({_al_u987_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [3]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,b_pad_gpio_porta_pad[3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u988_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [3]}),
    .q({open_n71502,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [3]}));  // ../RTL/gpio_ctrl.v(184)
  // ../RTL/gpio_apbif.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~A*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u989|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg6_b3  (
    .a({_al_u988_o,open_n71503}),
    .b({_al_u945_o,open_n71504}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [3],_al_u2490_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n61 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] ,\u_cmsdk_mcu/HWDATA [3]}),
    .mi({open_n71515,\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u989_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n195 }),
    .q({open_n71519,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/int_gpio_ls_sync [3]}));  // ../RTL/gpio_apbif.v(383)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u99 (
    .do({open_n71521,open_n71522,open_n71523,\u_cmsdk_mcu/p0_out [11]}),
    .ts(\u_cmsdk_mcu/p0_outen [11]),
    .opad(P0[11]));  // ../RTL/cmsdk_mcu_pin_mux.v(137)
  // ../RTL/gpio_apbif.v(363)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u990|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg5_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3],open_n71536}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [3],open_n71537}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,_al_u2492_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n58 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/HWDATA [3]}),
    .mi({open_n71548,\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u990_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n150 }),
    .q({open_n71552,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_int_polarity [3]}));  // ../RTL/gpio_apbif.v(363)
  // ../RTL/gpio_ctrl.v(248)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111001101011111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u991|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg3_b3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_intmask [3],open_n71553}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [3],open_n71554}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [3]}),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,_al_u3053_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u991_o,open_n71572}),
    .q({open_n71576,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [3]}));  // ../RTL/gpio_ctrl.v(248)
  // ../RTL/gpio_apbif.v(453)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u992|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg7_b3  (
    .b({_al_u990_o,_al_u992_o}),
    .c({_al_u991_o,_al_u994_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n68 ),
    .clk(XTAL1_wire),
    .d({_al_u566_o,_al_u989_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u992_o,open_n71595}),
    .q({open_n71599,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gpio0_prdata [3]}));  // ../RTL/gpio_apbif.v(453)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B*A))"),
    //.LUTF1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG0("(~D*~(~C*~B*A))"),
    //.LUTG1("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011111101),
    .INIT_LUTF1(16'b0000000010101100),
    .INIT_LUTG0(16'b0000000011111101),
    .INIT_LUTG1(16'b0000000010101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u993|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b3/B1_0 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }),
    .mi({open_n71603,\u_cmsdk_mcu/HADDR [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/sel0_b3/B1_0 ,_al_u994_o}),
    .q({open_n71618,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[6] }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/gpio_apbif.v(242)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(A*(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1010100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u996|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b2  (
    .a({_al_u470_o,open_n71619}),
    .b({b_pad_gpio_porta_pad[2],open_n71620}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2],_al_u2488_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2],\u_cmsdk_mcu/HWDATA [2]}),
    .mi({open_n71631,\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u996_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n238 }),
    .q({open_n71635,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [2]}));  // ../RTL/gpio_apbif.v(242)
  // ../RTL/gpio_apbif.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b1100100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u998|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg2_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [2],\u_cmsdk_mcu/HWDATA [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n63 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [2],_al_u3046_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n49 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_intr_ed_pm [2]}),
    .mi({open_n71646,\u_cmsdk_mcu/HWDATA [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_raw_intstatus [2],_al_u3047_o}),
    .q({open_n71650,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inten [2]}));  // ../RTL/gpio_apbif.v(303)
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u0|u1/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_0 ,1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_0 ,open_n71698}),
    .f({n0[0],open_n71718}),
    .fco(\u1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u10|u1/u9  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_9 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_9 }),
    .fci(\u1/c9 ),
    .f(n0[10:9]),
    .fco(\u1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u12|u1/u11  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_11 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_11 }),
    .fci(\u1/c11 ),
    .f(n0[12:11]),
    .fco(\u1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u13_al_u7271  (
    .a({open_n71767,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_13 }),
    .b({open_n71768,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_13 }),
    .fci(\u1/c13 ),
    .f({open_n71787,n0[13]}));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u2|u1/u1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_1 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_1 }),
    .fci(\u1/c1 ),
    .f(n0[2:1]),
    .fco(\u1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u4|u1/u3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_3 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_3 }),
    .fci(\u1/c3 ),
    .f(n0[4:3]),
    .fco(\u1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u6|u1/u5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_5 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_5 }),
    .fci(\u1/c5 ),
    .f(n0[6:5]),
    .fco(\u1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u8|u1/u7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_7 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_7 }),
    .fci(\u1/c7 ),
    .f(n0[8:7]),
    .fco(\u1/c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u0|u2/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_18 ,1'b0}),
    .b({n0[0],open_n71881}),
    .f({n1[0],open_n71901}),
    .fco(\u2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u10|u2/u9  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_28 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_27 }),
    .b(n0[10:9]),
    .fci(\u2/c9 ),
    .f(n1[10:9]),
    .fco(\u2/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u12|u2/u11  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_30 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_29 }),
    .b(n0[12:11]),
    .fci(\u2/c11 ),
    .f(n1[12:11]),
    .fco(\u2/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u13_al_u7272  (
    .a({open_n71950,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_31 }),
    .b({open_n71951,n0[13]}),
    .fci(\u2/c13 ),
    .f({open_n71970,n1[13]}));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u2|u2/u1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_20 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_19 }),
    .b(n0[2:1]),
    .fci(\u2/c1 ),
    .f(n1[2:1]),
    .fco(\u2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u4|u2/u3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_22 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_21 }),
    .b(n0[4:3]),
    .fci(\u2/c3 ),
    .f(n1[4:3]),
    .fco(\u2/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u6|u2/u5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_24 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_23 }),
    .b(n0[6:5]),
    .fci(\u2/c5 ),
    .f(n1[6:5]),
    .fco(\u2/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2/u0|u2/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2/u8|u2/u7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_26 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_25 }),
    .b(n0[8:7]),
    .fci(\u2/c7 ),
    .f(n1[8:7]),
    .fco(\u2/c9 ));
  EG_PHY_GCLK \u_M0clkpll/bufg_feedback  (
    .clki(\u_M0clkpll/clk0_buf ),
    .clko(XTAL1_wire));  // al_ip/M0clkpll.v(36)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(124),
    .CLKC0_DIV(125),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(1),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(3),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("ENABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u_M0clkpll/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(XTAL1_wire),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(XTAL1_pad),
    .reset(1'b0),
    .stdby(1'b0),
    .clkc({open_n72064,open_n72065,open_n72066,open_n72067,\u_M0clkpll/clk0_buf }));  // al_ip/M0clkpll.v(59)
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0004"),
    //.WID("0x0004"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_000  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_ram/n13 [8:0]),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa(\u_cmsdk_mcu/sram_hrdata [8:0]));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0005"),
    //.WID("0x0005"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_009  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_ram/n13 [17:9]),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa(\u_cmsdk_mcu/sram_hrdata [17:9]));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0006"),
    //.WID("0x0006"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_018  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_ram/n13 [26:18]),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa(\u_cmsdk_mcu/sram_hrdata [26:18]));
  // address_offset=0;data_offset=27;depth=1024;width=5;num_section=1;width_per_section=5;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0007"),
    //.WID("0x0007"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_ram/ram_memory0_1024x32_sub_000000_027  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia({open_n72152,open_n72153,open_n72154,open_n72155,5'b00000}),
    .dib({open_n72156,open_n72157,open_n72158,open_n72159,\u_cmsdk_mcu/u_ahb_ram/n13 [31:27]}),
    .web(\u_cmsdk_mcu/u_ahb_ram/n16 ),
    .doa({open_n72165,open_n72166,open_n72167,open_n72168,\u_cmsdk_mcu/sram_hrdata [31:27]}));
  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D)"),
    //.LUTF1("(~C*B*~(D*~A))"),
    //.LUTG0("(~D)"),
    //.LUTG1("(~C*B*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011111111),
    .INIT_LUTF1(16'b0000100000001100),
    .INIT_LUTG0(16'b0000000011111111),
    .INIT_LUTG1(16'b0000100000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_ahb_ram/reg0_b11|u_cmsdk_mcu/u_ahb_ram/reg0_b10  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uf9iu6 ,open_n72178}),
    .b({_al_u6286_o,open_n72179}),
    .c({_al_u6287_o,open_n72180}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .mi(\u_cmsdk_mcu/HADDR [11:10]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6288_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 }),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:10]));  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*~C))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000001000100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_ahb_ram/reg0_b12|u_cmsdk_mcu/u_ahb_ram/reg0_b4  (
    .a({open_n72198,_al_u6281_o}),
    .b({open_n72199,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bg9iu6 }),
    .c({\u_cmsdk_mcu/HADDR [12],\u_cmsdk_mcu/HADDR [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [13],\u_cmsdk_mcu/HADDR [4]}),
    .mi({\u_cmsdk_mcu/HADDR [12],\u_cmsdk_mcu/HADDR [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u4973_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uf9iu6 }),
    .q({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [12],\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [4]}));  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(~D*~C)))"),
    //.LUT1("(~D*(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010001001100),
    .INIT_LUT1(16'b0000000000111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_ahb_ram/reg0_b2|u_cmsdk_mcu/u_ahb_ram/reg0_b6  (
    .a({open_n72213,\u_cmsdk_mcu/HADDR [7]}),
    .b(\u_cmsdk_mcu/HADDR [7:6]),
    .c({\u_cmsdk_mcu/HADDR [2],\u_cmsdk_mcu/HADDR [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({_al_u5000_o,\u_cmsdk_mcu/HADDR [2]}),
    .mi({\u_cmsdk_mcu/HADDR [2],\u_cmsdk_mcu/HADDR [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6298_o,_al_u6287_o}),
    .q({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [2],\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [6]}));  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(C@B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~D*(C@B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000111100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_ahb_ram/reg0_b5|u_cmsdk_mcu/u_ahb_ram/reg0_b3  (
    .b({open_n72229,\u_cmsdk_mcu/HADDR [5]}),
    .c({\u_cmsdk_mcu/HADDR [5],\u_cmsdk_mcu/HADDR [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [8],_al_u5000_o}),
    .mi({\u_cmsdk_mcu/HADDR [5],\u_cmsdk_mcu/HADDR [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6284_o,_al_u6300_o}),
    .q({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [5],\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [3]}));  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~(B*A))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~D*~C*~(B*A))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000000000000111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_ahb_ram/reg0_b9|u_cmsdk_mcu/u_ahb_ram/reg0_b8  (
    .a({open_n72247,\u_cmsdk_mcu/HADDR [9]}),
    .b({\u_cmsdk_mcu/HADDR [8],\u_cmsdk_mcu/HADDR [8]}),
    .c({\u_cmsdk_mcu/HADDR [11],\u_cmsdk_mcu/HADDR [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [9],\u_cmsdk_mcu/HADDR [5]}),
    .mi(\u_cmsdk_mcu/HADDR [9:8]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6277_o,_al_u6279_o}),
    .q(\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [9:8]));  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*~D))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(~B*~(C*~D))"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011111100),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100110011111100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_ahb_ram/reg1_b0|u_cmsdk_mcu/u_ahb_ram/reg1_b16  (
    .b({open_n72267,\u_cmsdk_mcu/HSIZE [1]}),
    .c({\u_cmsdk_mcu/HADDR [1],\u_cmsdk_mcu/HADDR [1]}),
    .ce(\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [0],\u_cmsdk_mcu/HADDR [0]}),
    .f({\u_cmsdk_mcu/u_ahb_ram/n5 [0],open_n72285}),
    .q({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [16]}));  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*~D))"),
    //.LUTF1("~(~B*~(~C*~D))"),
    //.LUTG0("~(~B*~(C*~D))"),
    //.LUTG1("~(~B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011111100),
    .INIT_LUTF1(16'b1100110011001111),
    .INIT_LUTG0(16'b1100110011111100),
    .INIT_LUTG1(16'b1100110011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_ahb_ram/reg1_b10|u_cmsdk_mcu/u_ahb_ram/reg1_b24  (
    .b({\u_cmsdk_mcu/HSIZE [1],\u_cmsdk_mcu/HSIZE [1]}),
    .c({\u_cmsdk_mcu/HADDR [1],\u_cmsdk_mcu/HADDR [1]}),
    .ce(\u_cmsdk_mcu/u_ahb_ram/mux3_b0_sel_is_2_o ),
    .clk(XTAL1_wire),
    .d({_al_u5006_o,_al_u5006_o}),
    .q({\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [10],\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [24]}));  // ../RTL/AHB2MEM.v(51)
  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_ahb_ram/we_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b1  (
    .b({open_n72315,\u_cmsdk_mcu/u_cmsdk_mcu_system/sysrom_hsel }),
    .c({_al_u5003_o,\u_cmsdk_mcu/flash_hsel }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/sram_hsel ,_al_u5017_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({open_n72328,\u_cmsdk_mcu/sram_hsel }),
    .q({\u_cmsdk_mcu/u_ahb_ram/we ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [1]}));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0008"),
    //.WID("0x0008"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_000  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_rom/n13 [8:0]),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa(\u_cmsdk_mcu/flash_hrdata [8:0]));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0009"),
    //.WID("0x0009"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_009  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_rom/n13 [17:9]),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa(\u_cmsdk_mcu/flash_hrdata [17:9]));
  // address_offset=0;data_offset=18;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000A"),
    //.WID("0x000A"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_018  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia(9'b000000000),
    .dib(\u_cmsdk_mcu/u_ahb_rom/n13 [26:18]),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa(\u_cmsdk_mcu/flash_hrdata [26:18]));
  // address_offset=0;data_offset=27;depth=1024;width=5;num_section=1;width_per_section=5;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000B"),
    //.WID("0x000B"),
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("OFF"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("READBEFOREWRITE"))
    \u_cmsdk_mcu/u_ahb_rom/ram_memory0_1024x32_sub_000000_027  (
    .addra({\u_cmsdk_mcu/HADDR [11:2],3'b111}),
    .addrb({\u_cmsdk_mcu/u_ahb_ram/buf_hwaddr [11:2],3'b111}),
    .clka(XTAL1_wire),
    .clkb(XTAL1_wire),
    .dia({open_n72406,open_n72407,open_n72408,open_n72409,5'b00000}),
    .dib({open_n72410,open_n72411,open_n72412,open_n72413,\u_cmsdk_mcu/u_ahb_rom/n13 [31:27]}),
    .web(\u_cmsdk_mcu/u_ahb_rom/n16 ),
    .doa({open_n72419,open_n72420,open_n72421,open_n72422,\u_cmsdk_mcu/flash_hrdata [31:27]}));
  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  // ../RTL/AHB2MEM.v(51)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_ahb_rom/we_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg3_b0  (
    .c({_al_u5003_o,\u_cmsdk_mcu/u_ahb_ram/n5 [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/flash_hsel ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_ahb_rom/we ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_byte_strobe [0]}));  // ../RTL/cmsdk_mcu_sysctrl.v(147)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg_reg  (
    .clk(XTAL1_wire),
    .mi({open_n72469,1'b1}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .q({open_n72486,\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg }));  // ../RTL/cmsdk_mcu_clkctrl.v(108)
  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reg0_b1|u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reg0_b0  (
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [0],1'b1}),
    .sr(NRST_pad),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [1:0]));  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reg0_b2  (
    .clk(XTAL1_wire),
    .mi({open_n72530,\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [1]}),
    .sr(NRST_pad),
    .q({open_n72536,\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]}));  // ../RTL/cmsdk_mcu_clkctrl.v(86)
  // ../RTL/cortexm0ds_logic.v(17800)
  // ../RTL/cmsdk_ahb_to_iop.v(87)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~((D*C))*~(A)+B*(D*C)*~(A)+~(B)*(D*C)*A+B*(D*C)*A)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110010001000100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1110010001000100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/IOWRITE_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6_reg  (
    .a({open_n72537,_al_u5000_o}),
    .b({open_n72538,\u_cmsdk_mcu/HWRITE }),
    .c({\u_cmsdk_mcu/HWRITE ,_al_u5001_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HTRANS [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .mi({\u_cmsdk_mcu/HWRITE ,open_n72543}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u5003_o,open_n72555}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOWRITE ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }));  // ../RTL/cortexm0ds_logic.v(17800)
  // ../RTL/cortexm0ds_logic.v(17864)
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~A*~(D*C))"),
    //.LUTF1("(~D*(C@B))"),
    //.LUTG0("~(~B*~A*~(D*C))"),
    //.LUTG1("(~D*(C@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111011101110),
    .INIT_LUTF1(16'b0000000000111100),
    .INIT_LUTG0(16'b1111111011101110),
    .INIT_LUTG1(16'b0000000000111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b10|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6_reg  (
    .a({open_n72559,_al_u6295_o}),
    .b({\u_cmsdk_mcu/HADDR [10],_al_u6296_o}),
    .c({\u_cmsdk_mcu/HADDR [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5000_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }),
    .mi({\u_cmsdk_mcu/HADDR [10],open_n72564}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6296_o,open_n72576}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W5ypw6 }));  // ../RTL/cortexm0ds_logic.v(17864)
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~B*~(~D*~C)))"),
    //.LUTF1("(~A*~(~D*~(~C*B)))"),
    //.LUTG0("(~A*~(~B*~(~D*~C)))"),
    //.LUTG1("(~A*~(~D*~(~C*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010001000101),
    .INIT_LUTF1(16'b0101010100000100),
    .INIT_LUTG0(16'b0100010001000101),
    .INIT_LUTG1(16'b0101010100000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b11|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b4  (
    .a({_al_u6274_o,\u_cmsdk_mcu/HADDR [9]}),
    .b({_al_u6275_o,\u_cmsdk_mcu/HADDR [7]}),
    .c({\u_cmsdk_mcu/HADDR [8],\u_cmsdk_mcu/HADDR [4]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HADDR [11],\u_cmsdk_mcu/HADDR [3]}),
    .mi({\u_cmsdk_mcu/HADDR [11],\u_cmsdk_mcu/HADDR [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6276_o,_al_u6275_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b8|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b7  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8],\u_cmsdk_mcu/HADDR [8]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9],\u_cmsdk_mcu/HADDR [7]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7],\u_cmsdk_mcu/HADDR [10]}),
    .mi(\u_cmsdk_mcu/HADDR [8:7]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u580_o,_al_u6273_o}),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8:7]));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b1010101110101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b1  (
    .a({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [1]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [0],\u_cmsdk_mcu/p1_out [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/p1_out [0],\u_cmsdk_mcu/p1_out [1]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b1010101110101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b10|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b9  (
    .a(\u_cmsdk_mcu/HWDATA [10:9]),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 }),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [4:3]),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_out [10:9]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/p1_out [10:9]));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b1010101110101000),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b1010101110101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b11|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b8  (
    .a({\u_cmsdk_mcu/HWDATA [11],\u_cmsdk_mcu/HWDATA [8]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [11],\u_cmsdk_mcu/p1_out [8]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/p1_out [11],\u_cmsdk_mcu/p1_out [8]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b1010101110101000),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b1010101110101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b12|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b14  (
    .a({\u_cmsdk_mcu/HWDATA [12],\u_cmsdk_mcu/HWDATA [14]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [12],\u_cmsdk_mcu/p1_out [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/p1_out [12],\u_cmsdk_mcu/p1_out [14]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b1010101110101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b13|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b15  (
    .a({\u_cmsdk_mcu/HWDATA [13],\u_cmsdk_mcu/HWDATA [15]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write1 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n39 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [13],\u_cmsdk_mcu/p1_out [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/p1_out [13],\u_cmsdk_mcu/p1_out [15]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b1010101110101000),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b1010101110101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b2  (
    .a(\u_cmsdk_mcu/HWDATA [3:2]),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 }),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [5:4]),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/p1_out [3:2]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/p1_out [3:2]));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTF1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUTG1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101110101000),
    .INIT_LUTF1(16'b1010101110101000),
    .INIT_LUTG0(16'b1010101110101000),
    .INIT_LUTG1(16'b1010101110101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b4|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b6  (
    .a({\u_cmsdk_mcu/HWDATA [4],\u_cmsdk_mcu/HWDATA [6]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [4],\u_cmsdk_mcu/p1_out [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/p1_out [4],\u_cmsdk_mcu/p1_out [6]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(309)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b1010101110101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b5|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg1_b7  (
    .a({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [7]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_dout_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [9]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n34 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [5],\u_cmsdk_mcu/p1_out [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/p1_out [5],\u_cmsdk_mcu/p1_out [7]}));  // ../RTL/cmsdk_iop_gpio.v(309)
  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b15|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b15  (
    .a({open_n72766,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({open_n72767,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/p1_outen [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [15],\u_cmsdk_mcu/p1_out [15]}),
    .mi({open_n72772,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [15]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({open_n72784,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b15/B1_0 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [15]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b2  (
    .a({open_n72788,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({open_n72789,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/p1_outen [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [2],\u_cmsdk_mcu/p1_out [2]}),
    .mi({open_n72794,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({open_n72806,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b2/B1_0 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [2]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_iop_gpio.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000010000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011001000010000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg9_b6|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg0_b6  (
    .a({open_n72810,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}),
    .b({open_n72811,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [3]}),
    .c({\u_cmsdk_mcu/p1_outen [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/p1_out [6],\u_cmsdk_mcu/p1_out [6]}),
    .mi({open_n72816,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({open_n72828,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/mux0_b6/B1_0 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync1 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_in_sync2 [6]}));  // ../RTL/cmsdk_iop_gpio.v(252)
  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b5|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg0_b6  (
    .b({_al_u4977_o,_al_u4977_o}),
    .c({\u_cmsdk_mcu/HADDR [12],\u_cmsdk_mcu/HADDR [12]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/n11 ),
    .clk(XTAL1_wire),
    .d({_al_u4917_o,_al_u4917_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio0_hsel ,\u_cmsdk_mcu/u_cmsdk_mcu_system/gpio1_hsel }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [6]}));  // ../RTL/cmsdk_ahb_slave_mux.v(115)
  // ../RTL/gpio_apbif.v(343)
  // ../RTL/gpio_apbif.v(343)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg4_b2  (
    .c({_al_u2494_o,_al_u2494_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n55 ),
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3:2]),
    .mi(\u_cmsdk_mcu/HWDATA [3:2]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n105 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n103 }),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_inttype_level [3:2]));  // ../RTL/gpio_apbif.v(343)
  // ../RTL/gpio_apbif.v(242)
  // ../RTL/gpio_apbif.v(242)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b5|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/reg8_b3  (
    .c({_al_u2488_o,_al_u2488_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_apbif/n40 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [3]}),
    .mi({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n244 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n240 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_dr [3]}));  // ../RTL/gpio_apbif.v(242)
  // ../RTL/gpio_ctrl.v(203)
  // ../RTL/gpio_ctrl.v(192)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUT1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001000000010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b0  (
    .a({open_n72895,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [0]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3040_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [0]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [0]}));  // ../RTL/gpio_ctrl.v(203)
  // ../RTL/gpio_ctrl.v(203)
  // ../RTL/gpio_ctrl.v(192)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000000010),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b0011001000000010),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b1|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b1  (
    .a({open_n72910,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [1]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3075_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [1]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [1]}));  // ../RTL/gpio_ctrl.v(203)
  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(203)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000000010),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b0011001000000010),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b2  (
    .a({open_n72929,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3046_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [2]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [2]}));  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(203)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUT1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001000000010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b3  (
    .a({open_n72948,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3052_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [3]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [3]}));  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(203)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUT1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001000000010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b4|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b4  (
    .a({open_n72963,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [4]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3057_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [4]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [4]}));  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(203)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000000010),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b0011001000000010),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b5|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b5  (
    .a({open_n72978,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [5]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [5]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3062_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [5]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [5]}));  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(203)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000000010),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b0011001000000010),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b6|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b6  (
    .a({open_n72997,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [6]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3067_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [6]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [6]}));  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(192)
  // ../RTL/gpio_ctrl.v(203)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUT1("(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001000000010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg2_b7|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/reg1_b7  (
    .a({open_n73016,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/gpio_ext_porta_int [7]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_ls_sync }),
    .clk(1'b1),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/gpio_swporta_ddr [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_s1 [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3072_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ls_int_in [7]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/ed_int_d1 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_gpio_0$u_gpio_0/x_gpio_ctrl/int_pre_in [7]}));  // ../RTL/gpio_ctrl.v(192)
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [0],1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ,open_n73031}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .clk(XTAL1_wire),
    .mi({open_n73046,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [0],open_n73047}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c1 ),
    .q({open_n73050,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [2]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [2:1]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [2:1]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/u3_al_u7273  (
    .a({open_n73073,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_tick_cnt [3]}),
    .b({open_n73074,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add0/c3 ),
    .f({open_n73093,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n55 [3]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [0],1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_inc ,open_n73099}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [0],open_n73119}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [2:1]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [2:1]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/u3_al_u7274  (
    .a({open_n73146,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3]}),
    .b({open_n73147,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add1/c3 ),
    .f({open_n73166,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [3]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [0],1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ,open_n73172}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/BAUDTICK ),
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_2 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [0],open_n73187}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c1 ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_lpf [1:0]));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [2:1]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [2:1]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/u3_al_u7275  (
    .a({open_n73212,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [3]}),
    .b({open_n73213,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add2/c3 ),
    .f({open_n73232,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [3]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0],1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ,open_n73238}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .clk(XTAL1_wire),
    .mi(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [3:2]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [0],open_n73253}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c1 ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [2:1]));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2:1]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [2:1]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/u3_al_u7276  (
    .a({open_n73278,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]}),
    .b({open_n73279,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/add3/c3 ),
    .f({open_n73298,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [3]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_cin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [0],1'b1}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3],open_n73304}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [2:1]),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c1 ),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_cout|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_3  (
    .a({1'b0,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [3]}),
    .b({1'b1,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/lt0_c3 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n31 ,open_n73372}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    //.LUTF1("(~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    //.LUTG0("(A*~B*~C*D+~A*B*~C*D+~A*~B*C*D)"),
    //.LUTG1("(~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0001011000000000),
    .INIT_LUTF1(16'b1101010100000000),
    .INIT_LUTG0(16'b0001011000000000),
    .INIT_LUTG1(16'b1101010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b0_rom0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b3_rom0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [3]}));
  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("(A*~B*~C*D+~A*B*~C*D+A*~B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b1010011000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/mux4_b4_rom0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b4  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,open_n73402}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,_al_u478_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [4],open_n73415}),
    .q({open_n73419,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [4]}));  // ../RTL/cmsdk_apb_uart.v(303)
  // ../RTL/cmsdk_apb_uart.v(238)
  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b1  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable ,open_n73422}),
    .c({_al_u571_o,_al_u2488_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .clk(XTAL1_wire),
    .d({_al_u473_o,\u_cmsdk_mcu/HWDATA [1]}),
    .mi({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n236 }),
    .q({uart0_txen_pad,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]}));  // ../RTL/cmsdk_apb_uart.v(238)
  // ../RTL/cmsdk_apb_uart.v(238)
  // ../RTL/cmsdk_apb_uart.v(238)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B*D))"),
    //.LUT1("~(~C*~(B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011110000),
    .INIT_LUT1(16'b1111110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b5|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg0_b3  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable08 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [3]}),
    .mi({\u_cmsdk_mcu/HWDATA [5],\u_cmsdk_mcu/HWDATA [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n281 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n277 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [3]}));  // ../RTL/cmsdk_apb_uart.v(238)
  // ../RTL/cmsdk_apb_uart.v(583)
  // ../RTL/cmsdk_apb_uart.v(583)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("~(~D*~(C*B))"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("~(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b1111111111000000),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b1111111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b1|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b0  (
    .a({open_n73455,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 }),
    .b({_al_u364_o,_al_u364_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n88_lutinv }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ),
    .clk(XTAL1_wire),
    .d({_al_u560_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [0]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1:0]));  // ../RTL/cmsdk_apb_uart.v(583)
  // ../RTL/cmsdk_apb_uart.v(583)
  // ../RTL/cmsdk_apb_uart.v(583)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg10_b3  (
    .b({open_n73479,_al_u364_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n102 [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ),
    .clk(XTAL1_wire),
    .d({_al_u364_o,_al_u560_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [3]}));  // ../RTL/cmsdk_apb_uart.v(583)
  // ../RTL/cmsdk_apb_uart.v(603)
  // ../RTL/cmsdk_apb_uart.v(603)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b1|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg11_b2  (
    .b({open_n73503,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_buf_full }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxbuf_sample ),
    .clk(XTAL1_wire),
    .d({_al_u650_o,_al_u650_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n106 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_overrun }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_rx_buf [2]}));  // ../RTL/cmsdk_apb_uart.v(603)
  // ../RTL/cmsdk_apb_uart.v(614)
  // ../RTL/cmsdk_apb_uart.v(614)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*~A)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b4|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b3  (
    .a({open_n73517,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc }),
    .b({open_n73518,_al_u370_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n100 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state [1]}),
    .mi(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [5:4]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_update ,_al_u560_o}),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [4:3]));  // ../RTL/cmsdk_apb_uart.v(614)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg12_b5  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_state_inc ),
    .clk(XTAL1_wire),
    .mi({open_n73543,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({open_n73560,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_shift_buf [5]}));  // ../RTL/cmsdk_apb_uart.v(614)
  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(207)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*D))"),
    //.LUTF1("~(C*~D)"),
    //.LUTG0("~(~C*~(B*D))"),
    //.LUTG1("~(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011110000),
    .INIT_LUTF1(16'b1111111100001111),
    .INIT_LUTG0(16'b1111110011110000),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b6  (
    .b({open_n73563,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/reg_intclr_normal_write0 }),
    .c({_al_u637_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/new_masked_int [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({\u_cmsdk_mcu/HWDATA [0],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n50 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n283 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [6]}));  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(207)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b1|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b7  (
    .b({_al_u637_o,open_n73583}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_buf_full ,_al_u2488_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({\u_cmsdk_mcu/HWDATA [1],\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_overrun ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_iop_gpio/n248 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [7]}));  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(207)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b2  (
    .c({_al_u2484_o,_al_u2484_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [3:2]),
    .mi(\u_cmsdk_mcu/HWDATA [3:2]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n60 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n58 }),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [3:2]));  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(207)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b5|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg13_b4  (
    .c({_al_u2484_o,_al_u2484_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable00 ),
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [5:4]),
    .mi(\u_cmsdk_mcu/HWDATA [5:4]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n64 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n62 }),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [5:4]));  // ../RTL/cmsdk_apb_uart.v(207)
  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~C*B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000010000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b16|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b17  (
    .a({\u_cmsdk_mcu/HWDATA [30],open_n73643}),
    .b({\u_cmsdk_mcu/HWDATA [17],open_n73644}),
    .c({\u_cmsdk_mcu/HWDATA [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({_al_u3779_o,\u_cmsdk_mcu/HWDATA [17]}),
    .mi({\u_cmsdk_mcu/HWDATA [16],\u_cmsdk_mcu/HWDATA [17]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3780_o,_al_u3449_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [17]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cmsdk_apb_uart.v(247)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg1_b4  (
    .c({_al_u2482_o,_al_u2482_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/write_enable10 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/HWDATA [4]}),
    .mi({\u_cmsdk_mcu/HWDATA [3],\u_cmsdk_mcu/HWDATA [4]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n105 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n107 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [4]}));  // ../RTL/cmsdk_apb_uart.v(247)
  // ../RTL/cmsdk_apb_uart.v(303)
  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("~(D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("~(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b1100000011111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b1100000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b5  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .clk(XTAL1_wire),
    .d({_al_u494_o,_al_u475_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [5]}));  // ../RTL/cmsdk_apb_uart.v(303)
  // ../RTL/cmsdk_apb_uart.v(303)
  // ../RTL/cmsdk_apb_uart.v(303)
  EG_PHY_LSLICE #(
    //.LUTF0("((D*B)*~(C)*~(A)+(D*B)*C*~(A)+~((D*B))*C*A+(D*B)*C*A)"),
    //.LUTF1("~(~B*~((~D*~C))*~(A)+~B*(~D*~C)*~(A)+~(~B)*(~D*~C)*A+~B*(~D*~C)*A)"),
    //.LUTG0("((D*B)*~(C)*~(A)+(D*B)*C*~(A)+~((D*B))*C*A+(D*B)*C*A)"),
    //.LUTG1("~(~B*~((~D*~C))*~(A)+~B*(~D*~C)*~(A)+~(~B)*(~D*~C)*A+~B*(~D*~C)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110010010100000),
    .INIT_LUTF1(16'b1110111011100100),
    .INIT_LUTG0(16'b1110010010100000),
    .INIT_LUTG1(16'b1110111011100100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b1|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg2_b7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n25_lutinv }),
    .b({_al_u572_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n27_lutinv }),
    .c({_al_u573_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n26 [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_enable ),
    .clk(XTAL1_wire),
    .d({_al_u576_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/read_mux_byte0_reg [7]}));  // ../RTL/cmsdk_apb_uart.v(303)
  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b8  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [12]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [8]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [8]}));  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b10|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b7  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [11]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [7]}));  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b11|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b5  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [9]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [5]}));  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b12|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b4  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [16],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [8]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [12],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [4]}));  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b13|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b3  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [17],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [7]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [3]}));  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(341)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b14|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg3_b15  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_div [19]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [15]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n38 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [15]}));  // ../RTL/cmsdk_apb_uart.v(341)
  // ../RTL/cmsdk_apb_uart.v(358)
  // ../RTL/cmsdk_apb_uart.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("~(~C*D)"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("~(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b1111000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg4_b2  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n44 ),
    .clk(XTAL1_wire),
    .d({_al_u685_o,_al_u685_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2]}));  // ../RTL/cmsdk_apb_uart.v(358)
  // ../RTL/cmsdk_apb_uart.v(445)
  // ../RTL/cmsdk_apb_uart.v(445)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~A*~(D*~B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("~(~C*~A*~(D*~B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101111111010),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b1111101111111010),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg6_b1  (
    .a({open_n73870,_al_u1032_o}),
    .b({_al_u1035_o,_al_u1035_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n63 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state_update ),
    .clk(XTAL1_wire),
    .d({_al_u1032_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n67 [1]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_state [1]}));  // ../RTL/cmsdk_apb_uart.v(445)
  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(461)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b1|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b2  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [2]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .clk(XTAL1_wire),
    .d({_al_u637_o,_al_u637_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [2]}));  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(461)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b4  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [4]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [5]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .clk(XTAL1_wire),
    .d({_al_u637_o,_al_u637_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [4]}));  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(461)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b5|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b6  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [7]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .clk(XTAL1_wire),
    .d({_al_u637_o,_al_u637_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [6]}));  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(461)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b7|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg7_b0  (
    .b({open_n73955,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [0]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_tx_buf [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [1]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n74 ),
    .clk(XTAL1_wire),
    .d({_al_u637_o,_al_u637_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/tx_shift_buf [0]}));  // ../RTL/cmsdk_apb_uart.v(461)
  // ../RTL/cmsdk_apb_uart.v(535)
  // ../RTL/cmsdk_apb_uart.v(535)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b3  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [3]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ),
    .clk(XTAL1_wire),
    .d({_al_u388_o,_al_u388_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [3]}));  // ../RTL/cmsdk_apb_uart.v(535)
  // ../RTL/cmsdk_apb_uart.v(535)
  // ../RTL/cmsdk_apb_uart.v(535)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b1|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg9_b2  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n92 [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/update_rx_tick_cnt ),
    .clk(XTAL1_wire),
    .d({_al_u388_o,_al_u388_o}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rx_tick_cnt [2]}));  // ../RTL/cmsdk_apb_uart.v(535)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("CE"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("INV"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("SET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("ASYNC"),
    .TSMUX("1"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1_reg_IN  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_ctrl [1]),
    .ipad(uart0_rxd),
    .ipclk(XTAL1_wire),
    .rst(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .diq({open_n74028,open_n74029,open_n74030,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/rxd_sync_1 }));  // ../RTL/cmsdk_apb_uart.v(501)
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [0],1'b0}),
    .b({1'b1,open_n74033}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [0],open_n74053}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u10|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u9  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [10:9]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c9 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [10:9]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u12|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u11  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [12:11]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c11 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [12:11]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u14|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u13  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [14:13]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c13 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [14:13]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u15_al_u7277  (
    .a({open_n74124,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [15]}),
    .b({open_n74125,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c15 ),
    .f({open_n74144,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [15]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [2:1]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [2:1]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u4|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [4:3]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c3 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [4:3]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u6|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [6:5]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c5 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [6:5]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u8|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_i [8:7]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c7 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n37 [8:7]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub0/c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [0],1'b0}),
    .b({1'b1,open_n74238}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [0],open_n74258}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [2:1]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [2:1]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/u3_al_u7278  (
    .a({open_n74285,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/reg_baud_cntr_f [3]}),
    .b({open_n74286,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/sub1/c3 ),
    .f({open_n74305,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n43 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~D*~B*~C+~D*~B*C+~D*B*C)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/mux11_rom0|_al_u298  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1],open_n74313}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hreadyout }),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_slave_mux_sys_bus/reg_hsel [4]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hreadyout ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }));
  // ../RTL/cmsdk_ahb_to_apb.v(253)
  // ../RTL/cmsdk_ahb_to_apb.v(253)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTF1("(D*(C@B))"),
    //.LUTG0("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    //.LUTG1("(D*(C@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010111000111110),
    .INIT_LUTF1(16'b0011110000000000),
    .INIT_LUTG0(16'b0010111000111110),
    .INIT_LUTG1(16'b0011110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg2_b2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg2_b1  (
    .a({open_n74334,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 }),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [1:0]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2:1]),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/state_reg [2:1]));  // ../RTL/cmsdk_ahb_to_apb.v(253)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b1  (
    .b({open_n74359,\u_cmsdk_mcu/HADDR [3]}),
    .c({_al_u5009_o,\u_cmsdk_mcu/HADDR [2]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/apbsys_hsel ,_al_u6273_o}),
    .mi({\u_cmsdk_mcu/HADDR [2],\u_cmsdk_mcu/HADDR [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ,_al_u6274_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUTF1("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUTG0("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUTG1("(~A*~B*~C*D+A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001000000000),
    .INIT_LUTF1(16'b1010001100000000),
    .INIT_LUTG0(16'b1010001000000000),
    .INIT_LUTG1(16'b1010001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b2  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[2] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[3] }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] }),
    .mi(\u_cmsdk_mcu/HADDR [5:4]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/gen_apb_uart_0$u_apb_uart_0/n28 [7]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[4] }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~C*~B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b6|u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b8  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ,_al_u6277_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[9] ,_al_u6284_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] ,_al_u6285_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] ,\u_cmsdk_mcu/HADDR [10]}),
    .mi({\u_cmsdk_mcu/HADDR [8],\u_cmsdk_mcu/HADDR [10]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u465_o,_al_u6286_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[10] }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/u_ahb_to_apb/reg4_b9  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/n1 ),
    .clk(XTAL1_wire),
    .mi({open_n74425,\u_cmsdk_mcu/HADDR [11]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({open_n74431,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_apb_subsystem/PADDR[11] }));  // ../RTL/cmsdk_ahb_to_apb.v(153)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B*~C*D+~A*B*~C*D)"),
    //.LUT1("(~A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000010100000000),
    .INIT_LUT1(16'b1101010000000000),
    .MODE("LOGIC"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b0_rom0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/mux4_b1_rom0  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [0],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [1]}));
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B*~C*D+A*~B*C*D+A*B*C*D)"),
    //.LUT1("(A*~B*~C*D+~A*B*~C*D+A*~B*C*D+A*B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010001000000000),
    .INIT_LUT1(16'b1010011000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b3|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [2]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [4]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5]}),
    .mi({\u_cmsdk_mcu/HADDR [5],\u_cmsdk_mcu/HADDR [3]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [4],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/n19 [7]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [3]}));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b7|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b6  (
    .a({open_n74465,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [8]}),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [10:9]),
    .c(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [11:10]),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [11]}),
    .mi(\u_cmsdk_mcu/HADDR [9:8]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u496_o,_al_u4569_o}),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [9:8]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b9|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg0_b8  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/ahb_access ),
    .clk(XTAL1_wire),
    .mi(\u_cmsdk_mcu/HADDR [11:10]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cmsdk_mcu_sysctrl/reg_addr [11:10]));  // ../RTL/cmsdk_mcu_sysctrl.v(156)
  // ../RTL/cortexm0ds_logic.v(17778)
  // ../RTL/cortexm0ds_logic.v(17639)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A2spw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlvpw6_reg  (
    .a({open_n74510,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .b({open_n74511,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({open_n74512,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ,_al_u1155_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[19] }));  // ../RTL/cortexm0ds_logic.v(17778)
  // ../RTL/cortexm0ds_logic.v(18384)
  // ../RTL/cortexm0ds_logic.v(17185)
  EG_PHY_MSLICE #(
    //.LUT0("(C@D)"),
    //.LUT1("~(~B*~(C*~(D*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111110000),
    .INIT_LUT1(16'b1101110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ,open_n74527}),
    .b({_al_u3870_o,open_n74528}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 }),
    .mi({open_n74540,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsfax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({open_n74541,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A5ipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6 }));  // ../RTL/cortexm0ds_logic.v(18384)
  // ../RTL/cortexm0ds_logic.v(18904)
  // ../RTL/cortexm0ds_logic.v(18901)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acuax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xhuax6_reg  (
    .a({open_n74545,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({open_n74546,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({open_n74547,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc0pw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[7] }));  // ../RTL/cortexm0ds_logic.v(18904)
  // ../RTL/cortexm0ds_logic.v(17686)
  // ../RTL/cortexm0ds_logic.v(17630)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aurpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjtpw6_reg  (
    .a({open_n74562,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({open_n74563,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({open_n74564,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu2pw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[2] }));  // ../RTL/cortexm0ds_logic.v(17686)
  // ../RTL/cortexm0ds_logic.v(17648)
  // ../RTL/cortexm0ds_logic.v(19041)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,_al_u2508_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3fiu6 ,\u_cmsdk_mcu/HWDATA [14]}),
    .mi({\u_cmsdk_mcu/HWDATA [23],\u_cmsdk_mcu/HWDATA [14]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n82 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Auyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbspw6 }));  // ../RTL/cortexm0ds_logic.v(17648)
  // ../RTL/cortexm0ds_logic.v(19143)
  // ../RTL/cortexm0ds_logic.v(19149)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("~(C*D)"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6_reg  (
    .b({open_n74606,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5eiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u405_o,_al_u1883_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ,open_n74610}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R5eiu6 ,\u_cmsdk_mcu/HWDATA [0]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Avzax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zszax6 }));  // ../RTL/cortexm0ds_logic.v(19143)
  // ../RTL/cortexm0ds_logic.v(19849)
  // ../RTL/cortexm0ds_logic.v(19671)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,_al_u2476_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C0fiu6 ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({\u_cmsdk_mcu/HWDATA [30],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzeiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n246 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aw4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pz9bx6 }));  // ../RTL/cortexm0ds_logic.v(19849)
  // ../RTL/cortexm0ds_logic.v(19855)
  // ../RTL/cortexm0ds_logic.v(19575)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B*D))"),
    //.LUT1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011110000),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6_reg  (
    .b({open_n74644,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/reg_intclr_normal_write0 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/new_masked_int [6]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q0fiu6 ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ,\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n283 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Az3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R1abx6 }));  // ../RTL/cortexm0ds_logic.v(19855)
  // ../RTL/cortexm0ds_logic.v(17672)
  // ../RTL/cortexm0ds_logic.v(17638)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B0spw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z1tpw6_reg  (
    .a({open_n74658,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({open_n74659,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .c({open_n74660,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ,_al_u1197_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] }));  // ../RTL/cortexm0ds_logic.v(17672)
  // ../RTL/cortexm0ds_logic.v(20005)
  // ../RTL/cortexm0ds_logic.v(18897)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4uax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3fbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u789_o,_al_u786_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[22] }));  // ../RTL/cortexm0ds_logic.v(20005)
  // ../RTL/cortexm0ds_logic.v(18895)
  // ../RTL/cortexm0ds_logic.v(18898)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B6uax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D0uax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u833_o,_al_u861_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[2] }));  // ../RTL/cortexm0ds_logic.v(18895)
  // ../RTL/cortexm0ds_logic.v(18396)
  // ../RTL/cortexm0ds_logic.v(17331)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(D*~(C*B)))"),
    //.LUTF1("(D*~(~B*~(C*A)))"),
    //.LUTG0("~(~A*~(D*~(C*B)))"),
    //.LUTG1("(D*~(~B*~(C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111110101010),
    .INIT_LUTF1(16'b1110110000000000),
    .INIT_LUTG0(16'b1011111110101010),
    .INIT_LUTG1(16'b1110110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ,_al_u3320_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ,_al_u1253_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S63iu6_lutinv }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B7lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ryfax6 }));  // ../RTL/cortexm0ds_logic.v(18396)
  // ../RTL/cortexm0ds_logic.v(19792)
  // ../RTL/cortexm0ds_logic.v(18899)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B8uax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z78bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u852_o,_al_u738_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[15] }));  // ../RTL/cortexm0ds_logic.v(19792)
  // ../RTL/cortexm0ds_logic.v(17685)
  // ../RTL/cortexm0ds_logic.v(17232)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bbjpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xhtpw6_reg  (
    .a({open_n74751,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .b({open_n74752,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({open_n74753,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ,_al_u1579_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] }));  // ../RTL/cortexm0ds_logic.v(17685)
  // ../RTL/cortexm0ds_logic.v(18132)
  // ../RTL/cortexm0ds_logic.v(19972)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("~(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b1111001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6_reg  (
    .b({_al_u1718_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ro8ax6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,_al_u1695_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 }));  // ../RTL/cortexm0ds_logic.v(18132)
  // ../RTL/cortexm0ds_logic.v(19811)
  // ../RTL/cortexm0ds_logic.v(18100)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6_reg  (
    .b({_al_u1676_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1675_o,_al_u1675_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 }),
    .f({_al_u1826_o,_al_u1829_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bk7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q89bx6 }));  // ../RTL/cortexm0ds_logic.v(19811)
  // ../RTL/cortexm0ds_logic.v(18124)
  // ../RTL/cortexm0ds_logic.v(20019)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [8]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .f({_al_u5834_o,_al_u5822_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kl8ax6 }));  // ../RTL/cortexm0ds_logic.v(18124)
  // ../RTL/cortexm0ds_logic.v(20057)
  // ../RTL/cortexm0ds_logic.v(19581)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6_reg  (
    .a({\u_cmsdk_mcu/HWDATA [22],open_n74827}),
    .b({\u_cmsdk_mcu/HWDATA [23],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K66iu6 }),
    .c({_al_u2717_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y0gbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2721_o,\u_cmsdk_mcu/HWDATA [22]}),
    .mi(\u_cmsdk_mcu/HWDATA [23:22]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u3783_o,_al_u3481_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C14bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jdgbx6 }));  // ../RTL/cortexm0ds_logic.v(20057)
  // ../RTL/cortexm0ds_logic.v(17830)
  // ../RTL/cortexm0ds_logic.v(19766)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C27bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P2xpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u899_o,_al_u756_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[18] }));  // ../RTL/cortexm0ds_logic.v(17830)
  // ../RTL/cortexm0ds_logic.v(18905)
  // ../RTL/cortexm0ds_logic.v(18896)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2uax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wjuax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u858_o,_al_u798_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] }));  // ../RTL/cortexm0ds_logic.v(18905)
  // ../RTL/cortexm0ds_logic.v(17943)
  // ../RTL/cortexm0ds_logic.v(17858)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010111000111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0010111000111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6_reg  (
    .a({open_n74873,_al_u1253_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1689_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qj1qw6 }),
    .f({_al_u1690_o,_al_u1687_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gl1qw6 }));  // ../RTL/cortexm0ds_logic.v(17943)
  // ../RTL/cortexm0ds_logic.v(17457)
  // ../RTL/cortexm0ds_logic.v(19767)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C47bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ejnpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[31] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u898_o,_al_u849_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[31] }));  // ../RTL/cortexm0ds_logic.v(17457)
  // ../RTL/cortexm0ds_logic.v(19842)
  // ../RTL/cortexm0ds_logic.v(20043)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,_al_u2480_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzdiu6 ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({\u_cmsdk_mcu/HWDATA [22],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dv9iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n156 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv9bx6 }));  // ../RTL/cortexm0ds_logic.v(19842)
  // ../RTL/cortexm0ds_logic.v(17446)
  // ../RTL/cortexm0ds_logic.v(17808)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C5wpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gxmpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u744_o,_al_u869_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[3] }));  // ../RTL/cortexm0ds_logic.v(17446)
  // ../RTL/cortexm0ds_logic.v(17627)
  // ../RTL/cortexm0ds_logic.v(17809)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7wpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dorpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[7] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 }),
    .f({_al_u742_o,_al_u885_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[7] }));  // ../RTL/cortexm0ds_logic.v(17627)
  // ../RTL/cortexm0ds_logic.v(18971)
  // ../RTL/cortexm0ds_logic.v(19769)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C87bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxxax6_reg  (
    .a({open_n74963,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({open_n74964,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({open_n74965,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ,_al_u1228_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[30] }));  // ../RTL/cortexm0ds_logic.v(18971)
  // ../RTL/cortexm0ds_logic.v(18062)
  // ../RTL/cortexm0ds_logic.v(17810)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C9wpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P34qw6_reg  (
    .a({open_n74984,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({open_n74985,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({open_n74986,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ltmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C96pw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] }));  // ../RTL/cortexm0ds_logic.v(18062)
  // ../RTL/cortexm0ds_logic.v(18851)
  // ../RTL/cortexm0ds_logic.v(19770)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ca7bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qkrax6_reg  (
    .a({open_n75005,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({open_n75006,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .c({open_n75007,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ,_al_u1538_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[30] }));  // ../RTL/cortexm0ds_logic.v(18851)
  // ../RTL/cortexm0ds_logic.v(19793)
  // ../RTL/cortexm0ds_logic.v(17812)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cdwpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z98bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u741_o,_al_u736_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] }));  // ../RTL/cortexm0ds_logic.v(19793)
  // ../RTL/cortexm0ds_logic.v(17827)
  // ../RTL/cortexm0ds_logic.v(17775)
  EG_PHY_MSLICE #(
    //.LUT0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUT1("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010111000111111),
    .INIT_LUT1(16'b0010111000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6_reg  (
    .a({_al_u1253_o,_al_u1253_o}),
    .b({_al_u1676_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 }),
    .f({_al_u1710_o,_al_u1708_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cfvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gwwpw6 }));  // ../RTL/cortexm0ds_logic.v(17827)
  // ../RTL/cortexm0ds_logic.v(17641)
  // ../RTL/cortexm0ds_logic.v(19773)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cg7bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5spw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1630_o,_al_u1547_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] }));  // ../RTL/cortexm0ds_logic.v(17641)
  // ../RTL/cortexm0ds_logic.v(18758)
  // ../RTL/cortexm0ds_logic.v(18740)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cglax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfmax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2246_o,_al_u2165_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u2247_o,_al_u2166_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[17] }));  // ../RTL/cortexm0ds_logic.v(18758)
  // ../RTL/cortexm0ds_logic.v(18906)
  // ../RTL/cortexm0ds_logic.v(19774)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ci7bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wluax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u1085_o,_al_u1211_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[26] }));  // ../RTL/cortexm0ds_logic.v(18906)
  // ../RTL/cortexm0ds_logic.v(17534)
  // ../RTL/cortexm0ds_logic.v(19775)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ck7bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9ppw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u897_o,_al_u850_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] }));  // ../RTL/cortexm0ds_logic.v(17534)
  // ../RTL/cortexm0ds_logic.v(18933)
  // ../RTL/cortexm0ds_logic.v(19777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Co7bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M3wax6_reg  (
    .a({open_n75124,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({open_n75125,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({open_n75126,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ,_al_u796_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[24] }));  // ../RTL/cortexm0ds_logic.v(18933)
  // ../RTL/cortexm0ds_logic.v(18964)
  // ../RTL/cortexm0ds_logic.v(17711)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*B))"),
    //.LUT1("~(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011111111),
    .INIT_LUT1(16'b1100000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8eiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [23],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [7]}),
    .clk(XTAL1_wire),
    .d({_al_u2312_o,_al_u2345_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 }));  // ../RTL/cortexm0ds_logic.v(18964)
  // ../RTL/cortexm0ds_logic.v(19953)
  // ../RTL/cortexm0ds_logic.v(18045)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [9]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .f({_al_u5832_o,_al_u5820_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cq3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlcbx6 }));  // ../RTL/cortexm0ds_logic.v(19953)
  // ../RTL/cortexm0ds_logic.v(17527)
  // ../RTL/cortexm0ds_logic.v(17628)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cqrpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ovopw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[29] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u1955_o,_al_u2423_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[29] }));  // ../RTL/cortexm0ds_logic.v(17527)
  // ../RTL/cortexm0ds_logic.v(19760)
  // ../RTL/cortexm0ds_logic.v(19761)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs6bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dq6bx6_reg  (
    .a({open_n75202,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({open_n75203,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztmiu6 ,_al_u846_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[8] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[9] }));  // ../RTL/cortexm0ds_logic.v(19760)
  // ../RTL/cortexm0ds_logic.v(17326)
  // ../RTL/cortexm0ds_logic.v(17492)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("~(B*A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b1111011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6_reg  (
    .a({_al_u1829_o,_al_u1823_o}),
    .b({_al_u1830_o,_al_u1824_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 }));  // ../RTL/cortexm0ds_logic.v(17326)
  // ../RTL/cortexm0ds_logic.v(19719)
  // ../RTL/cortexm0ds_logic.v(19749)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D46bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nk5bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u778_o,_al_u1208_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] }));  // ../RTL/cortexm0ds_logic.v(19719)
  // ../RTL/cortexm0ds_logic.v(19716)
  // ../RTL/cortexm0ds_logic.v(19750)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D66bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe5bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u774_o,_al_u840_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[6] }));  // ../RTL/cortexm0ds_logic.v(19716)
  // ../RTL/cortexm0ds_logic.v(19718)
  // ../RTL/cortexm0ds_logic.v(19751)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D86bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ni5bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[24] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u761_o,_al_u797_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] }));  // ../RTL/cortexm0ds_logic.v(19718)
  // ../RTL/cortexm0ds_logic.v(18951)
  // ../RTL/cortexm0ds_logic.v(19752)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Da6bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J3xax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u754_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5pow6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[4] }));  // ../RTL/cortexm0ds_logic.v(18951)
  // ../RTL/cortexm0ds_logic.v(18950)
  // ../RTL/cortexm0ds_logic.v(19753)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dc6bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K1xax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u749_o,_al_u864_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[2] }));  // ../RTL/cortexm0ds_logic.v(18950)
  // ../RTL/cortexm0ds_logic.v(18972)
  // ../RTL/cortexm0ds_logic.v(19754)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/De6bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzxax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u1244_o,_al_u1234_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[31] }));  // ../RTL/cortexm0ds_logic.v(18972)
  // ../RTL/cortexm0ds_logic.v(18225)
  // ../RTL/cortexm0ds_logic.v(18224)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L03qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ud4iu6 ,open_n75347}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cf7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dfbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgbax6 }));  // ../RTL/cortexm0ds_logic.v(18225)
  // ../RTL/cortexm0ds_logic.v(19757)
  // ../RTL/cortexm0ds_logic.v(19755)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg6bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dk6bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u732_o,_al_u718_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[12] }));  // ../RTL/cortexm0ds_logic.v(19757)
  // ../RTL/cortexm0ds_logic.v(19736)
  // ../RTL/cortexm0ds_logic.v(19756)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di6bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy5bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[25] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u725_o,_al_u802_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] }));  // ../RTL/cortexm0ds_logic.v(19736)
  // ../RTL/cortexm0ds_logic.v(17311)
  // ../RTL/cortexm0ds_logic.v(19961)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ,open_n75384}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wt3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ,_al_u1723_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2cbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Stkpw6 }),
    .f({_al_u367_o,_al_u1724_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvkpw6 }));  // ../RTL/cortexm0ds_logic.v(17311)
  // ../RTL/cortexm0ds_logic.v(17520)
  // ../RTL/cortexm0ds_logic.v(17795)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("~(B*A*~(D*C))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("~(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b1111011101110111),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b1111011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ir6ow6 }),
    .b({_al_u1652_o,_al_u1654_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P91ju6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G81ju6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jckax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wkipw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dzvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Shopw6 }));  // ../RTL/cortexm0ds_logic.v(17520)
  // ../RTL/cortexm0ds_logic.v(17453)
  // ../RTL/cortexm0ds_logic.v(17448)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1npw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ebnpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u816_o,_al_u720_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] }));  // ../RTL/cortexm0ds_logic.v(17453)
  // ../RTL/cortexm0ds_logic.v(20104)
  // ../RTL/cortexm0ds_logic.v(18565)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(~D*A))"),
    //.LUTF1("~(~(~C*B)*~(D*A))"),
    //.LUTG0("(~(~C*B)*~(~D*A))"),
    //.LUTG1("~(~(~C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001101010001),
    .INIT_LUTF1(16'b1010111000001100),
    .INIT_LUTG0(16'b1111001101010001),
    .INIT_LUTG1(16'b1010111000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6_reg  (
    .a({_al_u6746_o,_al_u6746_o}),
    .b({_al_u6743_o,_al_u6743_o}),
    .c({_al_u4530_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sn7iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E6iax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W8hbx6 }));  // ../RTL/cortexm0ds_logic.v(20104)
  // ../RTL/cortexm0ds_logic.v(19931)
  // ../RTL/cortexm0ds_logic.v(18089)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("~(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b1111001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6_reg  (
    .b({_al_u1701_o,_al_u1706_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z67ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdbbx6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufbbx6 }));  // ../RTL/cortexm0ds_logic.v(19931)
  // ../RTL/cortexm0ds_logic.v(17660)
  // ../RTL/cortexm0ds_logic.v(17452)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E9npw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ynspw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u1109_o,_al_u1187_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[24] }));  // ../RTL/cortexm0ds_logic.v(17660)
  // ../RTL/cortexm0ds_logic.v(18355)
  // ../RTL/cortexm0ds_logic.v(18343)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yc7iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rc7iu6 ,_al_u2040_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eafax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hdfax6 }));  // ../RTL/cortexm0ds_logic.v(18355)
  // ../RTL/cortexm0ds_logic.v(18881)
  // ../RTL/cortexm0ds_logic.v(18883)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0000000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ectax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F8tax6_reg  (
    .b({open_n75516,_al_u2423_o}),
    .c({open_n75517,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Csmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ,_al_u2424_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[25] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] }));  // ../RTL/cortexm0ds_logic.v(18881)
  // ../RTL/cortexm0ds_logic.v(17929)
  // ../RTL/cortexm0ds_logic.v(17454)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ednpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tu0qw6_reg  (
    .a({open_n75532,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .b({open_n75533,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jkniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[8] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Numiu6 ,_al_u882_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[8] }));  // ../RTL/cortexm0ds_logic.v(17929)
  // ../RTL/cortexm0ds_logic.v(17225)
  // ../RTL/cortexm0ds_logic.v(17456)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehnpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uwipw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1232_o,_al_u1091_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[31] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[4] }));  // ../RTL/cortexm0ds_logic.v(17225)
  // ../RTL/cortexm0ds_logic.v(18073)
  // ../RTL/cortexm0ds_logic.v(17462)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hqgiu6 ,\u_cmsdk_mcu/HWDATA [23]}),
    .mi({\u_cmsdk_mcu/HWDATA [31],\u_cmsdk_mcu/HWDATA [23]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Aqgiu6 ,_al_u3487_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Elnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 }));  // ../RTL/cortexm0ds_logic.v(18073)
  // ../RTL/cortexm0ds_logic.v(17777)
  // ../RTL/cortexm0ds_logic.v(17626)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emrpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjvpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({_al_u886_o,_al_u759_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] }));  // ../RTL/cortexm0ds_logic.v(17777)
  // ../RTL/cortexm0ds_logic.v(18868)
  // ../RTL/cortexm0ds_logic.v(18888)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Emtax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Misax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[2] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u2168_o,_al_u1913_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[2] }));  // ../RTL/cortexm0ds_logic.v(18868)
  // ../RTL/cortexm0ds_logic.v(18870)
  // ../RTL/cortexm0ds_logic.v(18891)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Estax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmsax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[23] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .f({_al_u2100_o,_al_u2246_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[23] }));  // ../RTL/cortexm0ds_logic.v(18870)
  // ../RTL/cortexm0ds_logic.v(18949)
  // ../RTL/cortexm0ds_logic.v(17950)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ez1qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lzwax6_reg  (
    .a({open_n75633,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({open_n75634,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Miniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jsmiu6 ,_al_u880_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[8] }));  // ../RTL/cortexm0ds_logic.v(18949)
  // ../RTL/cortexm0ds_logic.v(20173)
  // ../RTL/cortexm0ds_logic.v(17949)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fx1qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjibx6_reg  (
    .a({open_n75653,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({open_n75654,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[28] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Finiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qsmiu6 ,_al_u1221_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[28] }));  // ../RTL/cortexm0ds_logic.v(20173)
  // ../RTL/cortexm0ds_logic.v(17445)
  // ../RTL/cortexm0ds_logic.v(17447)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzmpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gvmpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({_al_u873_o,_al_u831_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[30] }));  // ../RTL/cortexm0ds_logic.v(17445)
  // ../RTL/cortexm0ds_logic.v(20132)
  // ../RTL/cortexm0ds_logic.v(19059)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6_reg  (
    .b({open_n75693,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fpgiu6 ,_al_u1935_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4eiu6 ,open_n75704}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P3fiu6 ,\u_cmsdk_mcu/HWDATA [4]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G0zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqhbx6 }));  // ../RTL/cortexm0ds_logic.v(20132)
  // ../RTL/cortexm0ds_logic.v(17384)
  // ../RTL/cortexm0ds_logic.v(17382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(C*D)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6_reg  (
    .b({open_n75710,_al_u3324_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U5yhu6 ,_al_u1676_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u530_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U03iu6 ,_al_u3325_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 }));  // ../RTL/cortexm0ds_logic.v(17384)
  // ../RTL/cortexm0ds_logic.v(17932)
  // ../RTL/cortexm0ds_logic.v(17948)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gv1qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q01qw6_reg  (
    .a({open_n75729,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({open_n75730,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Etmiu6 ,_al_u1602_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[8] }));  // ../RTL/cortexm0ds_logic.v(17932)
  // ../RTL/cortexm0ds_logic.v(17826)
  // ../RTL/cortexm0ds_logic.v(19763)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*D))"),
    //.LUT1("~(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001100110011),
    .INIT_LUT1(16'b1111001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6_reg  (
    .b({_al_u1692_o,_al_u1708_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bu6bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kswpw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Puwpw6 }));  // ../RTL/cortexm0ds_logic.v(17826)
  // ../RTL/cortexm0ds_logic.v(17661)
  // ../RTL/cortexm0ds_logic.v(18068)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gx6ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ypspw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u1178_o,_al_u1186_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[24] }));  // ../RTL/cortexm0ds_logic.v(17661)
  // ../RTL/cortexm0ds_logic.v(18320)
  // ../RTL/cortexm0ds_logic.v(18323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(~C*~B)*~(~D*~A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(~C*~B)*~(~D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111110010101000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111110010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6_reg  (
    .a({_al_u4035_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({_al_u4121_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lk9ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .f({_al_u5799_o,_al_u6754_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gzeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rteax6 }));  // ../RTL/cortexm0ds_logic.v(18320)
  // ../RTL/cortexm0ds_logic.v(20107)
  // ../RTL/cortexm0ds_logic.v(17325)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(D*C*~B))"),
    //.LUT1("~(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111010101010101),
    .INIT_LUT1(16'b1100000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6_reg  (
    .a({open_n75806,_al_u5836_o}),
    .b({_al_u5053_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .clk(XTAL1_wire),
    .d({_al_u5668_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H3lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 }));  // ../RTL/cortexm0ds_logic.v(20107)
  // ../RTL/cortexm0ds_logic.v(18965)
  // ../RTL/cortexm0ds_logic.v(17776)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(D*~(C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6_reg  (
    .b({_al_u2217_o,open_n75828}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F6eiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2210_o,\u_cmsdk_mcu/HWDATA [2]}),
    .f({\u_cmsdk_mcu/HWDATA [19],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3eiu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vlxax6 }));  // ../RTL/cortexm0ds_logic.v(18965)
  // ../RTL/cortexm0ds_logic.v(17774)
  // ../RTL/cortexm0ds_logic.v(17816)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*D))"),
    //.LUTF1("~(D*~(C*B))"),
    //.LUTG0("~(B*~(C*D))"),
    //.LUTG1("~(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100110011),
    .INIT_LUTF1(16'b1100000011111111),
    .INIT_LUTG0(16'b1111001100110011),
    .INIT_LUTG1(16'b1100000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,_al_u1710_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gbvpw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1704_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldvpw6 }));  // ../RTL/cortexm0ds_logic.v(17774)
  // ../RTL/cortexm0ds_logic.v(20260)
  // ../RTL/cortexm0ds_logic.v(18237)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(D*~(C*B)))"),
    //.LUT1("(C*~(B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111101010101),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6_reg  (
    .a({open_n75870,_al_u4452_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Scbiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmbax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lmkbx6 }));  // ../RTL/cortexm0ds_logic.v(20260)
  // ../RTL/cortexm0ds_logic.v(17930)
  // ../RTL/cortexm0ds_logic.v(17850)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hmxpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sw0qw6_reg  (
    .a({open_n75889,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .b({open_n75890,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ckniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gumiu6 ,_al_u1190_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[8] }));  // ../RTL/cortexm0ds_logic.v(17930)
  // ../RTL/cortexm0ds_logic.v(17154)
  // ../RTL/cortexm0ds_logic.v(17160)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6_reg  (
    .clk(SWCLKTCK_pad),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6 ,1'b1}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Evhpw6 }));  // ../RTL/cortexm0ds_logic.v(17154)
  // ../RTL/cortexm0ds_logic.v(17566)
  // ../RTL/cortexm0ds_logic.v(17490)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+~(D)*B*~(C)+D*B*~(C)+D*B*C)"),
    //.LUT1("~(B*~(C*~(D*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111100001100),
    .INIT_LUT1(16'b0111001111110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Di1iu6 ,open_n75933}),
    .b({_al_u3882_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Li7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 }));  // ../RTL/cortexm0ds_logic.v(17566)
  // ../RTL/cortexm0ds_logic.v(17831)
  // ../RTL/cortexm0ds_logic.v(17548)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I1qpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4xpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u1166_o,_al_u1151_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[18] }));  // ../RTL/cortexm0ds_logic.v(17831)
  // ../RTL/cortexm0ds_logic.v(17673)
  // ../RTL/cortexm0ds_logic.v(17549)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3qpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z3tpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u771_o,_al_u801_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] }));  // ../RTL/cortexm0ds_logic.v(17673)
  // ../RTL/cortexm0ds_logic.v(17704)
  // ../RTL/cortexm0ds_logic.v(17550)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5qpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y9upw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u723_o,_al_u747_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[17] }));  // ../RTL/cortexm0ds_logic.v(17704)
  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cortexm0ds_logic.v(18956)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("~(~D*~A*~(~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b1111111110101011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/u_ahb_to_gpio/reg0_b2  (
    .a({_al_u6295_o,open_n75994}),
    .b({_al_u5000_o,\u_cmsdk_mcu/HADDR [3]}),
    .c({\u_cmsdk_mcu/HADDR [4],\u_cmsdk_mcu/HADDR [2]}),
    .clk(XTAL1_wire),
    .d({_al_u6302_o,\u_cmsdk_mcu/HADDR [4]}),
    .mi({open_n76006,\u_cmsdk_mcu/HADDR [2]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({open_n76007,_al_u6281_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I5xax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_0/IOADDR [2]}));  // ../RTL/cmsdk_ahb_to_iop.v(78)
  // ../RTL/cortexm0ds_logic.v(17688)
  // ../RTL/cortexm0ds_logic.v(17551)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I7qpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Untpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({_al_u1097_o,_al_u1064_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[2] }));  // ../RTL/cortexm0ds_logic.v(17688)
  // ../RTL/cortexm0ds_logic.v(18274)
  // ../RTL/cortexm0ds_logic.v(18282)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(~C*~B)*~(~D*~A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(~C*~B)*~(~D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111110010101000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111110010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6_reg  (
    .a({_al_u4136_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u4225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eudax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S54iu6 }),
    .f({_al_u5712_o,_al_u6696_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iddax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lycax6 }));  // ../RTL/cortexm0ds_logic.v(18274)
  // ../RTL/cortexm0ds_logic.v(20183)
  // ../RTL/cortexm0ds_logic.v(18169)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wskhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Orkhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xajbx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 }),
    .f({_al_u5485_o,_al_u5239_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Im9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3jbx6 }));  // ../RTL/cortexm0ds_logic.v(20183)
  // ../RTL/cortexm0ds_logic.v(17547)
  // ../RTL/cortexm0ds_logic.v(17546)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ixppw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Izppw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u1217_o,_al_u1241_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] }));  // ../RTL/cortexm0ds_logic.v(17547)
  // ../RTL/cortexm0ds_logic.v(19945)
  // ../RTL/cortexm0ds_logic.v(18398)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("~(~B*~(D*C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b1101110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ,_al_u3320_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 }),
    .mi({open_n76089,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J4cbx6 }),
    .f({open_n76091,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J0gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A6cbx6 }));  // ../RTL/cortexm0ds_logic.v(19945)
  // ../RTL/cortexm0ds_logic.v(19951)
  // ../RTL/cortexm0ds_logic.v(18302)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6_reg  (
    .a({_al_u4096_o,open_n76095}),
    .b({_al_u4219_o,_al_u5095_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .f({_al_u5761_o,_al_u5096_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thcbx6 }));  // ../RTL/cortexm0ds_logic.v(19951)
  // ../RTL/cortexm0ds_logic.v(18187)
  // ../RTL/cortexm0ds_logic.v(20184)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(~C*B)*~(D@A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(~C*B)*~(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1010001001010001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1010001001010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I9ihu6 ,open_n76114}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A8ihu6 ,open_n76115}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C2ypw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ,open_n76119}),
    .f({_al_u5577_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J5jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yjaax6 }));  // ../RTL/cortexm0ds_logic.v(18187)
  // ../RTL/cortexm0ds_logic.v(17857)
  // ../RTL/cortexm0ds_logic.v(19974)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*B))"),
    //.LUTF1("~(D*~(C*B))"),
    //.LUTG0("~(D*~(C*B))"),
    //.LUTG1("~(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011111111),
    .INIT_LUTF1(16'b1100000011111111),
    .INIT_LUTG0(16'b1100000011111111),
    .INIT_LUTG1(16'b1100000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cydbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gyxpw6 }),
    .clk(SWCLKTCK_pad),
    .d({_al_u1713_o,_al_u1690_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L0ypw6 }));  // ../RTL/cortexm0ds_logic.v(17857)
  // ../RTL/cortexm0ds_logic.v(17526)
  // ../RTL/cortexm0ds_logic.v(17779)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jnvpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Otopw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u2211_o,_al_u1514_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] }));  // ../RTL/cortexm0ds_logic.v(17526)
  // ../RTL/cortexm0ds_logic.v(17663)
  // ../RTL/cortexm0ds_logic.v(17780)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jpvpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ytspw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[24] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u2215_o,_al_u2437_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[24] }));  // ../RTL/cortexm0ds_logic.v(17663)
  // ../RTL/cortexm0ds_logic.v(17676)
  // ../RTL/cortexm0ds_logic.v(17781)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jrvpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z9tpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u1156_o,_al_u1198_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[25] }));  // ../RTL/cortexm0ds_logic.v(17676)
  // ../RTL/cortexm0ds_logic.v(17840)
  // ../RTL/cortexm0ds_logic.v(17787)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*C)*~(~B*A))"),
    //.LUT1("~(~(D*C)*~(~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001000100010),
    .INIT_LUT1(16'b1111001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6_reg  (
    .a({_al_u5706_o,_al_u5706_o}),
    .b({_al_u5810_o,_al_u5814_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvvpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pexpw6 }));  // ../RTL/cortexm0ds_logic.v(17840)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kfoax6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kdkiu6 ),
    .clk(XTAL1_wire),
    .mi({open_n76235,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 }),
    .q({open_n76253,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[23] }));  // ../RTL/cortexm0ds_logic.v(18794)
  // ../RTL/cortexm0ds_logic.v(18871)
  // ../RTL/cortexm0ds_logic.v(18873)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kssax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kosax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hhqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[30] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy2pw6 ,_al_u2264_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[30] }));  // ../RTL/cortexm0ds_logic.v(18871)
  // ../RTL/cortexm0ds_logic.v(17560)
  // ../RTL/cortexm0ds_logic.v(17396)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~B*D)"),
    //.LUT1("(C*~(~B*~(~D*A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111111111),
    .INIT_LUT1(16'b1100000011100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6_reg  (
    .a({_al_u3869_o,open_n76272}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pmlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tezhu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfqpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({_al_u3870_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jq3iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 }));  // ../RTL/cortexm0ds_logic.v(17560)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6_reg  (
    .clk(SWCLKTCK_pad),
    .mi({open_n76298,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hwhpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/reset_sync_reg [2]),
    .q({open_n76315,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 }));  // ../RTL/cortexm0ds_logic.v(17166)
  // ../RTL/cortexm0ds_logic.v(17617)
  // ../RTL/cortexm0ds_logic.v(18718)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6_reg  (
    .a({open_n76316,_al_u4534_o}),
    .b({_al_u6746_o,_al_u4535_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/A25iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u6744_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L4lax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hgrpw6 }));  // ../RTL/cortexm0ds_logic.v(17617)
  // ../RTL/cortexm0ds_logic.v(19071)
  // ../RTL/cortexm0ds_logic.v(19083)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 ,open_n76339}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G2fiu6 ,open_n76340}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I45bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S1fiu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6689_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L1fiu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L8zax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H4zax6 }));  // ../RTL/cortexm0ds_logic.v(19071)
  // ../RTL/cortexm0ds_logic.v(19861)
  // ../RTL/cortexm0ds_logic.v(20063)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(C*D)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6_reg  (
    .b({open_n76360,\u_cmsdk_mcu/sram_hrdata [6]}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 ,\u_cmsdk_mcu/u_ahb_ram/hwdata_mask [0]}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ,\u_cmsdk_mcu/HWDATA [6]}),
    .mi({\u_cmsdk_mcu/HWDATA [22],\u_cmsdk_mcu/HWDATA [6]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ,\u_cmsdk_mcu/u_ahb_ram/n13 [6]}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3abx6 }));  // ../RTL/cortexm0ds_logic.v(19861)
  // ../RTL/cortexm0ds_logic.v(18930)
  // ../RTL/cortexm0ds_logic.v(18939)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lfwax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pxvax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[5] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u779_o,_al_u876_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] }));  // ../RTL/cortexm0ds_logic.v(18930)
  // ../RTL/cortexm0ds_logic.v(18255)
  // ../RTL/cortexm0ds_logic.v(19815)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111101001100),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6_reg  (
    .a({_al_u4066_o,_al_u4111_o}),
    .b({_al_u4141_o,_al_u4141_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yybax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .f({_al_u5740_o,_al_u5744_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J8cax6 }));  // ../RTL/cortexm0ds_logic.v(18255)
  // ../RTL/cortexm0ds_logic.v(18927)
  // ../RTL/cortexm0ds_logic.v(18940)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lhwax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rrvax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[31] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .f({_al_u1161_o,_al_u1235_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[31] }));  // ../RTL/cortexm0ds_logic.v(18927)
  // ../RTL/cortexm0ds_logic.v(18090)
  // ../RTL/cortexm0ds_logic.v(19889)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTF1("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTG1("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001111101111),
    .INIT_LUTF1(16'b0010111000111111),
    .INIT_LUTG0(16'b0010001111101111),
    .INIT_LUTG1(16'b0010111000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6_reg  (
    .a({_al_u1253_o,_al_u1253_o}),
    .b({_al_u1676_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E97ax6 }),
    .f({_al_u1699_o,_al_u1701_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Liabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Va7ax6 }));  // ../RTL/cortexm0ds_logic.v(18090)
  // ../RTL/cortexm0ds_logic.v(17664)
  // ../RTL/cortexm0ds_logic.v(17539)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljppw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yvspw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u1168_o,_al_u1184_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[24] }));  // ../RTL/cortexm0ds_logic.v(17664)
  // ../RTL/cortexm0ds_logic.v(18935)
  // ../RTL/cortexm0ds_logic.v(18941)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljwax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M7wax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u762_o,_al_u815_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] }));  // ../RTL/cortexm0ds_logic.v(18935)
  // ../RTL/cortexm0ds_logic.v(17834)
  // ../RTL/cortexm0ds_logic.v(17540)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llppw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Paxpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[18] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 }),
    .f({_al_u1160_o,_al_u1148_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[18] }));  // ../RTL/cortexm0ds_logic.v(17834)
  // ../RTL/cortexm0ds_logic.v(18947)
  // ../RTL/cortexm0ds_logic.v(18942)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Llwax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lvwax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[12] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 }),
    .f({_al_u755_o,_al_u719_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] }));  // ../RTL/cortexm0ds_logic.v(18947)
  // ../RTL/cortexm0ds_logic.v(17533)
  // ../RTL/cortexm0ds_logic.v(17541)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lnppw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N7ppw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[30] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 }),
    .f({_al_u1107_o,_al_u1227_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[30] }));  // ../RTL/cortexm0ds_logic.v(17533)
  // ../RTL/cortexm0ds_logic.v(17536)
  // ../RTL/cortexm0ds_logic.v(17542)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lpppw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mdppw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[5] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1096_o,_al_u1103_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[5] }));  // ../RTL/cortexm0ds_logic.v(17536)
  // ../RTL/cortexm0ds_logic.v(20008)
  // ../RTL/cortexm0ds_logic.v(18934)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M5wax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9fbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wk5pw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ml6pw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] }));  // ../RTL/cortexm0ds_logic.v(20008)
  // ../RTL/cortexm0ds_logic.v(17939)
  // ../RTL/cortexm0ds_logic.v(17936)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b1100000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6_reg  (
    .b({_al_u5053_o,_al_u5820_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pl4iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5258_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M81qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 }));  // ../RTL/cortexm0ds_logic.v(17939)
  // ../RTL/cortexm0ds_logic.v(19599)
  // ../RTL/cortexm0ds_logic.v(19611)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 ,open_n76577}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1fiu6 ,open_n76578}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2fiu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6687_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mb4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74bx6 }));  // ../RTL/cortexm0ds_logic.v(19599)
  // ../RTL/cortexm0ds_logic.v(18411)
  // ../RTL/cortexm0ds_logic.v(18281)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010000101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6_reg  (
    .a({_al_u4197_o,open_n76596}),
    .b({_al_u4231_o,open_n76597}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2rpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ,open_n76608}),
    .f({_al_u5719_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yogax6 }));  // ../RTL/cortexm0ds_logic.v(18411)
  // ../RTL/cortexm0ds_logic.v(18938)
  // ../RTL/cortexm0ds_logic.v(18937)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mbwax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ldwax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V6now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wanow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E8now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u768_o,_al_u804_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[25] }));  // ../RTL/cortexm0ds_logic.v(18938)
  // ../RTL/cortexm0ds_logic.v(20100)
  // ../RTL/cortexm0ds_logic.v(18313)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6_reg  (
    .a({_al_u4091_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({_al_u4191_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zt1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wxgbx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .f({_al_u5802_o,_al_u6797_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mgeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1hbx6 }));  // ../RTL/cortexm0ds_logic.v(20100)
  // ../RTL/cortexm0ds_logic.v(17940)
  // ../RTL/cortexm0ds_logic.v(17941)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b1111001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6_reg  (
    .b({_al_u5246_o,_al_u5818_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5053_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mh1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 }));  // ../RTL/cortexm0ds_logic.v(17940)
  // ../RTL/cortexm0ds_logic.v(17675)
  // ../RTL/cortexm0ds_logic.v(17429)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mjmpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z7tpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2441_o,_al_u2255_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u2442_o,_al_u2256_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] }));  // ../RTL/cortexm0ds_logic.v(17675)
  // ../RTL/cortexm0ds_logic.v(17449)
  // ../RTL/cortexm0ds_logic.v(18712)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0lax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E3npw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Panow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[29] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({_al_u711_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rt4pw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[29] }));  // ../RTL/cortexm0ds_logic.v(17449)
  // ../RTL/cortexm0ds_logic.v(18779)
  // ../RTL/cortexm0ds_logic.v(18787)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N1oax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nlnax6_reg  (
    .a({open_n76704,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({open_n76705,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gq4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r12_o[29] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dhniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ,_al_u1531_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[29] }));  // ../RTL/cortexm0ds_logic.v(18779)
  // ../RTL/cortexm0ds_logic.v(18294)
  // ../RTL/cortexm0ds_logic.v(18301)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("((D@B)*(C@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0001001001001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6_reg  (
    .a({_al_u4066_o,_al_u1916_o}),
    .b({_al_u4121_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 }),
    .f({_al_u5770_o,_al_u2201_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3eax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kqdax6 }));  // ../RTL/cortexm0ds_logic.v(18294)
  // ../RTL/cortexm0ds_logic.v(18178)
  // ../RTL/cortexm0ds_logic.v(18400)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(C*B)*~(~D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111100010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mzihu6 ,open_n76734}),
    .b({_al_u5598_o,open_n76735}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lm1iu6 ,open_n76746}),
    .f({_al_u5604_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T94iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N4gax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2aax6 }));  // ../RTL/cortexm0ds_logic.v(18178)
  // ../RTL/cortexm0ds_logic.v(19814)
  // ../RTL/cortexm0ds_logic.v(18182)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*B)*~(~D*A))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001101010001),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C4ihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M1ihu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jraax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 }),
    .f({_al_u5581_o,_al_u5539_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Naaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pe9bx6 }));  // ../RTL/cortexm0ds_logic.v(19814)
  // ../RTL/cortexm0ds_logic.v(20105)
  // ../RTL/cortexm0ds_logic.v(18406)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhlhu6 ,open_n76765}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gglhu6 ,open_n76766}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nv3qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 ,open_n76770}),
    .f({_al_u5497_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M94iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nfgax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wahbx6 }));  // ../RTL/cortexm0ds_logic.v(20105)
  // ../RTL/cortexm0ds_logic.v(18782)
  // ../RTL/cortexm0ds_logic.v(18777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nhnax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nrnax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .f({_al_u2449_o,_al_u2219_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[20] }));  // ../RTL/cortexm0ds_logic.v(18782)
  // ../RTL/cortexm0ds_logic.v(20000)
  // ../RTL/cortexm0ds_logic.v(19720)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nm5bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ttebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jjwow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pdyow6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[22] }));  // ../RTL/cortexm0ds_logic.v(20000)
  // ../RTL/cortexm0ds_logic.v(18181)
  // ../RTL/cortexm0ds_logic.v(19891)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oeihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmihu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Clihu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cndbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .f({_al_u5561_o,_al_u5564_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q8aax6 }));  // ../RTL/cortexm0ds_logic.v(18181)
  // ../RTL/cortexm0ds_logic.v(19892)
  // ../RTL/cortexm0ds_logic.v(20015)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010000101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6_reg  (
    .a({_al_u4086_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u4131_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Esabx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P74iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L54iu6 }),
    .f({_al_u5753_o,_al_u6720_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nnfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Koabx6 }));  // ../RTL/cortexm0ds_logic.v(19892)
  // ../RTL/cortexm0ds_logic.v(18299)
  // ../RTL/cortexm0ds_logic.v(18293)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("((D@B)*(C@A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("((D@B)*(C@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001001001000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001001001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6_reg  (
    .a({_al_u4071_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u4111_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 }),
    .f({_al_u5776_o,_al_u5223_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nodax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzdax6 }));  // ../RTL/cortexm0ds_logic.v(18299)
  // ../RTL/cortexm0ds_logic.v(19764)
  // ../RTL/cortexm0ds_logic.v(18133)
  EG_PHY_MSLICE #(
    //.LUT0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001111101111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6_reg  (
    .a({open_n76868,_al_u1253_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1694_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wq8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gw6bx6 }),
    .f({_al_u1695_o,_al_u1692_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xx6bx6 }));  // ../RTL/cortexm0ds_logic.v(19764)
  // ../RTL/cortexm0ds_logic.v(19810)
  // ../RTL/cortexm0ds_logic.v(19983)
  EG_PHY_MSLICE #(
    //.LUT0("~((C*~B)*~(D)*~(A)+(C*~B)*D*~(A)+~((C*~B))*D*A+(C*~B)*D*A)"),
    //.LUT1("(~D*~C*~(~B*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010111101111),
    .INIT_LUT1(16'b0000000000001101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ufebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [1]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 }),
    .f({_al_u4953_o,_al_u5836_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nwdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B79bx6 }));  // ../RTL/cortexm0ds_logic.v(19810)
  // ../RTL/cortexm0ds_logic.v(17674)
  // ../RTL/cortexm0ds_logic.v(17530)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O1ppw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z5tpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[25] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u1402_o,_al_u1498_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[25] }));  // ../RTL/cortexm0ds_logic.v(17674)
  // ../RTL/cortexm0ds_logic.v(17430)
  // ../RTL/cortexm0ds_logic.v(18861)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O4sax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mlmpw6_reg  (
    .a({open_n76915,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2283_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[27] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .f({_al_u2284_o,_al_u2445_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[27] }));  // ../RTL/cortexm0ds_logic.v(17430)
  // ../RTL/cortexm0ds_logic.v(17707)
  // ../RTL/cortexm0ds_logic.v(17532)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O5ppw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfupw6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[4] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] }));  // ../RTL/cortexm0ds_logic.v(17707)
  // ../RTL/cortexm0ds_logic.v(18772)
  // ../RTL/cortexm0ds_logic.v(18775)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Odnax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R7nax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jo4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Drkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1610_o,_al_u1586_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[3] }));  // ../RTL/cortexm0ds_logic.v(18772)
  // ../RTL/cortexm0ds_logic.v(17643)
  // ../RTL/cortexm0ds_logic.v(18856)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ourax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9spw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[6] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u2233_o,_al_u1950_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[6] }));  // ../RTL/cortexm0ds_logic.v(17643)
  // ../RTL/cortexm0ds_logic.v(19980)
  // ../RTL/cortexm0ds_logic.v(18321)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6_reg  (
    .a({_al_u4076_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dw1iu6 }),
    .b({_al_u4111_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ar1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fjdbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J44iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .f({_al_u5804_o,_al_u5179_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oveax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqdbx6 }));  // ../RTL/cortexm0ds_logic.v(19980)
  // ../RTL/cortexm0ds_logic.v(18849)
  // ../RTL/cortexm0ds_logic.v(18857)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Owrax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rgrax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[4] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u2223_o,_al_u1932_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[4] }));  // ../RTL/cortexm0ds_logic.v(18849)
  // ../RTL/cortexm0ds_logic.v(20002)
  // ../RTL/cortexm0ds_logic.v(17529)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ozopw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Txebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ds4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rs4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r8_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u1458_o,_al_u1474_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[22] }));  // ../RTL/cortexm0ds_logic.v(20002)
  // ../RTL/cortexm0ds_logic.v(17694)
  // ../RTL/cortexm0ds_logic.v(17833)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P8xpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xztpw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ljqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2202_o,_al_u2449_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u2203_o,_al_u2450_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[26] }));  // ../RTL/cortexm0ds_logic.v(17694)
  // ../RTL/cortexm0ds_logic.v(17493)
  // ../RTL/cortexm0ds_logic.v(18025)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1681_o,_al_u1675_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 }),
    .f({_al_u1683_o,_al_u1681_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P93qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3opw6 }));  // ../RTL/cortexm0ds_logic.v(17493)
  // ../RTL/cortexm0ds_logic.v(20185)
  // ../RTL/cortexm0ds_logic.v(18260)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~C*~B)*~(~D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111110010101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6_reg  (
    .a({_al_u4225_o,open_n77072}),
    .b({_al_u4237_o,open_n77073}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 }),
    .f({_al_u5739_o,_al_u1979_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Phcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F7jbx6 }));  // ../RTL/cortexm0ds_logic.v(20185)
  // ../RTL/cortexm0ds_logic.v(18360)
  // ../RTL/cortexm0ds_logic.v(18359)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(~(A)*~(B)*~(D)+A*B*D))"),
    //.LUTF1("~(~C*~B*~D)"),
    //.LUTG0("(C*(~(A)*~(B)*~(D)+A*B*D))"),
    //.LUTG1("~(~C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000010000),
    .INIT_LUTF1(16'b1111111111111100),
    .INIT_LUTG0(16'b1000000000010000),
    .INIT_LUTG1(16'b1111111111111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6_reg  (
    .a({open_n77088,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzlpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z73qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D2opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zgfax6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pifax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Okfax6 }));  // ../RTL/cortexm0ds_logic.v(18360)
  // ../RTL/cortexm0ds_logic.v(18222)
  // ../RTL/cortexm0ds_logic.v(20255)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jf7iu6 ,open_n77111}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 ,open_n77112}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tikbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sg7iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 }),
    .f({_al_u5656_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lg7iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pkkbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lbbax6 }));  // ../RTL/cortexm0ds_logic.v(18222)
  // ../RTL/cortexm0ds_logic.v(17695)
  // ../RTL/cortexm0ds_logic.v(17883)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Plypw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1upw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .f({_al_u765_o,_al_u807_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[26] }));  // ../RTL/cortexm0ds_logic.v(17695)
  // ../RTL/cortexm0ds_logic.v(20097)
  // ../RTL/cortexm0ds_logic.v(18174)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W9lhu6 ,open_n77145}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjkhu6 ,open_n77146}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ,open_n77150}),
    .f({_al_u5504_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pv9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvgbx6 }));  // ../RTL/cortexm0ds_logic.v(20097)
  // ../RTL/cortexm0ds_logic.v(17287)
  // ../RTL/cortexm0ds_logic.v(18710)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pwkax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T3kpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nq4ju6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wr4ju6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ls9pw6 ,_al_u1594_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[5] }));  // ../RTL/cortexm0ds_logic.v(17287)
  // ../RTL/cortexm0ds_logic.v(17908)
  // ../RTL/cortexm0ds_logic.v(20181)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pzibx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xozpw6_reg  (
    .b({_al_u1551_o,_al_u1586_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 }),
    .f({_al_u1552_o,_al_u1587_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[1] }));  // ../RTL/cortexm0ds_logic.v(17908)
  // ../RTL/cortexm0ds_logic.v(20103)
  // ../RTL/cortexm0ds_logic.v(19968)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("(~D*~C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6_reg  (
    .a({_al_u4549_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oa4iu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bvfbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [6]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W74iu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fs6iu6 ,_al_u5826_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H7hbx6 }));  // ../RTL/cortexm0ds_logic.v(20103)
  // ../RTL/cortexm0ds_logic.v(20081)
  // ../RTL/cortexm0ds_logic.v(19623)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*B*~(~C*A))"),
    //.LUT1("(~D*~(B*~(~C*A)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011000100),
    .INIT_LUT1(16'b0000000000111011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F5uow6 }),
    .b({_al_u6388_o,_al_u6388_o}),
    .c({_al_u6389_o,_al_u6389_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N2fiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 }),
    .mi({\u_cmsdk_mcu/HWDATA [30],\u_cmsdk_mcu/HWDATA [22]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6399_o,_al_u6400_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qf4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rlgbx6 }));  // ../RTL/cortexm0ds_logic.v(20081)
  // ../RTL/cortexm0ds_logic.v(19982)
  // ../RTL/cortexm0ds_logic.v(19952)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6_reg  (
    .a({_al_u4076_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .b({_al_u4096_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zodbx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .f({_al_u5725_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hcuiu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qudbx6 }));  // ../RTL/cortexm0ds_logic.v(19982)
  // ../RTL/cortexm0ds_logic.v(18999)
  // ../RTL/cortexm0ds_logic.v(19011)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 ,open_n77247}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ,_al_u2484_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X0fiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6527_o,\u_cmsdk_mcu/HWDATA [7]}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fsdiu6 ,\u_cmsdk_mcu/HWDATA [7]}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({_al_u6528_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n68 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qjyax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mfyax6 }));  // ../RTL/cortexm0ds_logic.v(18999)
  // ../RTL/cortexm0ds_logic.v(17662)
  // ../RTL/cortexm0ds_logic.v(17522)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qlopw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yrspw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u2264_o,_al_u2433_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K39iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zvkiu6 }),
    .f({_al_u2265_o,_al_u2434_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[24] }));  // ../RTL/cortexm0ds_logic.v(17662)
  // ../RTL/cortexm0ds_logic.v(18410)
  // ../RTL/cortexm0ds_logic.v(18292)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~(~C*~B)*~(~D*~A))"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~(~C*~B)*~(~D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b1111110010101000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b1111110010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6_reg  (
    .a({_al_u4184_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 }),
    .b({_al_u4197_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D84iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F94iu6 }),
    .f({_al_u5774_o,_al_u922_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qmdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bngax6 }));  // ../RTL/cortexm0ds_logic.v(18410)
  // ../RTL/cortexm0ds_logic.v(17521)
  // ../RTL/cortexm0ds_logic.v(17524)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qpopw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rjopw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1919_o,_al_u1928_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1920_o,_al_u1929_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[4] }));  // ../RTL/cortexm0ds_logic.v(17521)
  // ../RTL/cortexm0ds_logic.v(17881)
  // ../RTL/cortexm0ds_logic.v(18709)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qukax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhypw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qiqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ofkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jy2pw6 ,_al_u1964_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tx8iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 }),
    .f({_al_u1875_o,_al_u1965_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[0] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r9_o[1] }));  // ../RTL/cortexm0ds_logic.v(17881)
  // ../RTL/cortexm0ds_logic.v(18924)
  // ../RTL/cortexm0ds_logic.v(18929)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qvvax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Slvax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jgkiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ef8iu6 }),
    .f({_al_u1077_o,_al_u1089_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[4] }));  // ../RTL/cortexm0ds_logic.v(18924)
  // ../RTL/cortexm0ds_logic.v(17581)
  // ../RTL/cortexm0ds_logic.v(18390)
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    //.LUT1("(~(D@C)*~(B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000001111),
    .INIT_LUT1(16'b0111000000000111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6_reg  (
    .a({_al_u1255_o,open_n77357}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Krlpw6 ,open_n77358}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qufax6 ,open_n77370}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S63iu6_lutinv ,open_n77371}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 }));  // ../RTL/cortexm0ds_logic.v(17581)
  // ../RTL/cortexm0ds_logic.v(17390)
  // ../RTL/cortexm0ds_logic.v(17484)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(~C*B*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001111111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qynpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6_reg  (
    .b({open_n77377,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Golpw6 }),
    .c({_al_u368_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vplpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u367_o,_al_u3259_o}),
    .mi({open_n77381,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L5lpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({open_n77393,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W13iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P13iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oulpw6 }));  // ../RTL/cortexm0ds_logic.v(17390)
  // ../RTL/cortexm0ds_logic.v(18145)
  // ../RTL/cortexm0ds_logic.v(18157)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111111111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6_reg  (
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4rpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 ,open_n77404}),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bs4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R19ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 }));  // ../RTL/cortexm0ds_logic.v(18145)
  // ../RTL/cortexm0ds_logic.v(17723)
  // ../RTL/cortexm0ds_logic.v(18981)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6_reg  (
    .a({_al_u6295_o,_al_u6295_o}),
    .b({_al_u6300_o,_al_u6298_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eh6iu6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R9yax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ztupw6 }));  // ../RTL/cortexm0ds_logic.v(17723)
  // ../RTL/cortexm0ds_logic.v(17595)
  // ../RTL/cortexm0ds_logic.v(17971)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTF1("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTG0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG1("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010111000111111),
    .INIT_LUTF1(16'b0010001111101111),
    .INIT_LUTG0(16'b0010111000111111),
    .INIT_LUTG1(16'b0010001111101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6_reg  (
    .a({_al_u1253_o,_al_u1253_o}),
    .b({_al_u1676_o,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S02iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay1iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ra2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yzqpw6 }));  // ../RTL/cortexm0ds_logic.v(17595)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkpw6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Afkiu6 ),
    .clk(XTAL1_wire),
    .mi({open_n77473,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .q({open_n77480,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r11_o[21] }));  // ../RTL/cortexm0ds_logic.v(17297)
  // ../RTL/cortexm0ds_logic.v(18921)
  // ../RTL/cortexm0ds_logic.v(20172)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rhibx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vfvax6_reg  (
    .a({open_n77481,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({open_n77482,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Khniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[9] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vjniu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K3niu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xsmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y1xow6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[28] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[9] }));  // ../RTL/cortexm0ds_logic.v(18921)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("A7"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("INV"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("SET"),
    .IOTYPE("LVCMOS25"),
    .MODE("BI"),
    .SRMODE("ASYNC"),
    .TSMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6_reg_IN  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tw2iu6 ),
    .do({open_n77501,open_n77502,open_n77503,\u_cmsdk_mcu/dbg_swdo }),
    .ipclk(SWCLKTCK_pad),
    .rst(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .ts(\u_cmsdk_mcu/dbg_swdo_en ),
    .diq({open_n77509,open_n77510,open_n77511,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rilpw6 }),
    .bpad(SWDIOTMS));  // ../RTL/cmsdk_mcu.v(167)
  // ../RTL/cortexm0ds_logic.v(19795)
  // ../RTL/cortexm0ds_logic.v(18925)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rnvax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zd8bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rdkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vx9iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y50pw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[15] }));  // ../RTL/cortexm0ds_logic.v(19795)
  // ../RTL/cortexm0ds_logic.v(19799)
  // ../RTL/cortexm0ds_logic.v(20178)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rtibx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zl8bx6_reg  (
    .b({_al_u1519_o,_al_u1415_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gfniu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1520_o,_al_u1416_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[13] }));  // ../RTL/cortexm0ds_logic.v(19799)
  // ../RTL/cortexm0ds_logic.v(18275)
  // ../RTL/cortexm0ds_logic.v(18272)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(~C*~B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0101010010101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6_reg  (
    .a({_al_u4066_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .b({_al_u4126_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vr1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bwdax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E54iu6 }),
    .f({_al_u5711_o,_al_u6733_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rucax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 }));  // ../RTL/cortexm0ds_logic.v(18275)
  // ../RTL/cortexm0ds_logic.v(18257)
  // ../RTL/cortexm0ds_logic.v(19806)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6_reg  (
    .a({_al_u4116_o,open_n77561}),
    .b({_al_u4121_o,open_n77562}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cs1iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q44iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gk4iu6 }),
    .f({_al_u5757_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rz8bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bccax6 }));  // ../RTL/cortexm0ds_logic.v(18257)
  // ../RTL/cortexm0ds_logic.v(19885)
  // ../RTL/cortexm0ds_logic.v(17410)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6_reg  (
    .c({_al_u2482_o,_al_u2482_o}),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B3fiu6 ),
    .clk(XTAL1_wire),
    .d(\u_cmsdk_mcu/HWDATA [7:6]),
    .mi(\u_cmsdk_mcu/HWDATA [7:6]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n113 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_ahb_gpio_1/u_iop_gpio/n111 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3mpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcabx6 }));  // ../RTL/cortexm0ds_logic.v(19885)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S3nax6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mekiu6 ),
    .clk(XTAL1_wire),
    .mi({open_n77616,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D39iu6 }),
    .q({open_n77623,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r14_o[31] }));  // ../RTL/cortexm0ds_logic.v(18770)
  // ../RTL/cortexm0ds_logic.v(20006)
  // ../RTL/cortexm0ds_logic.v(18116)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S58ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T5fbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X7now6_lutinv }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N9now6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ddkiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u729_o,_al_u783_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] }));  // ../RTL/cortexm0ds_logic.v(20006)
  // ../RTL/cortexm0ds_logic.v(20012)
  // ../RTL/cortexm0ds_logic.v(18118)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S98ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Thfbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ep4ju6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ydkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u1408_o,_al_u1472_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u1409_o,_al_u1473_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_psp_o[20] }));  // ../RTL/cortexm0ds_logic.v(20012)
  // ../RTL/cortexm0ds_logic.v(17545)
  // ../RTL/cortexm0ds_logic.v(17880)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sfypw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jvppw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[5] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1142_o,_al_u1100_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[5] }));  // ../RTL/cortexm0ds_logic.v(17545)
  // ../RTL/cortexm0ds_logic.v(17909)
  // ../RTL/cortexm0ds_logic.v(17926)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/So0qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wqzpw6_reg  (
    .b({_al_u1602_o,_al_u1594_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X6niu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rkkiu6 }),
    .f({_al_u1603_o,_al_u1595_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[3] }));  // ../RTL/cortexm0ds_logic.v(17909)
  // ../RTL/cortexm0ds_logic.v(19395)
  // ../RTL/cortexm0ds_logic.v(19551)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*B))"),
    //.LUT1("(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000001010000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6_reg  (
    .a({_al_u3874_o,_al_u3874_o}),
    .b({\u_cmsdk_mcu/HWDATA [8],\u_cmsdk_mcu/HWDATA [1]}),
    .c({_al_u3935_o,_al_u3932_o}),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kwfiu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sq3bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y72bx6 }));  // ../RTL/cortexm0ds_logic.v(19395)
  // ../RTL/cortexm0ds_logic.v(19997)
  // ../RTL/cortexm0ds_logic.v(18112)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sx7ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tnebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dmqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u1121_o,_al_u1174_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[22] }));  // ../RTL/cortexm0ds_logic.v(19997)
  // ../RTL/cortexm0ds_logic.v(19998)
  // ../RTL/cortexm0ds_logic.v(18113)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sz7ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tpebx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[22] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mx8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 }),
    .f({_al_u1118_o,_al_u1175_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[22] }));  // ../RTL/cortexm0ds_logic.v(19998)
  // ../RTL/cortexm0ds_logic.v(17172)
  // ../RTL/cortexm0ds_logic.v(17178)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*~(B*~(D*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ehqpw6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq ,\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F42iu6 ,_al_u3319_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T0ipw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nyhpw6 }));  // ../RTL/cortexm0ds_logic.v(17172)
  // ../RTL/cortexm0ds_logic.v(17910)
  // ../RTL/cortexm0ds_logic.v(17917)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T60qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vszpw6_reg  (
    .b({_al_u1463_o,_al_u1543_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1464_o,_al_u1544_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[4] }));  // ../RTL/cortexm0ds_logic.v(17910)
  // ../RTL/cortexm0ds_logic.v(17925)
  // ../RTL/cortexm0ds_logic.v(17919)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ta0qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tm0qw6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,_al_u1618_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({_al_u1448_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hymiu6 }),
    .f({_al_u1449_o,_al_u1619_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[8] }));  // ../RTL/cortexm0ds_logic.v(17925)
  // ../RTL/cortexm0ds_logic.v(18423)
  // ../RTL/cortexm0ds_logic.v(18030)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~A*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~A*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0001010100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0001010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf1iu6 ,open_n77796}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nmfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gpqpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V34iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/H34iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5816_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/M24iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tb3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 }));  // ../RTL/cortexm0ds_logic.v(18423)
  // ../RTL/cortexm0ds_logic.v(17922)
  // ../RTL/cortexm0ds_logic.v(17920)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc0qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tg0qw6_reg  (
    .b({_al_u1439_o,_al_u1423_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n1552 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lp4ju6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 }),
    .f({_al_u1440_o,_al_u1424_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_msp_o[14] }));  // ../RTL/cortexm0ds_logic.v(17922)
  // ../RTL/cortexm0ds_logic.v(18163)
  // ../RTL/cortexm0ds_logic.v(19813)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q4lhu6 ,open_n77830}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qnkhu6 ,open_n77831}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kw1iu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xi4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .f({_al_u5477_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tc9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ab9ax6 }));  // ../RTL/cortexm0ds_logic.v(18163)
  // ../RTL/cortexm0ds_logic.v(18271)
  // ../RTL/cortexm0ds_logic.v(20188)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(~D*~A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(~D*~A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100101010),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011111100101010),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6_reg  (
    .a({_al_u4071_o,_al_u4071_o}),
    .b({_al_u4237_o,_al_u4126_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I0dax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Md7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ym4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .f({_al_u5718_o,_al_u5713_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tcjbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uscax6 }));  // ../RTL/cortexm0ds_logic.v(18271)
  // ../RTL/cortexm0ds_logic.v(17691)
  // ../RTL/cortexm0ds_logic.v(17879)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tdypw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xttpw6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fzkiu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[26] }));  // ../RTL/cortexm0ds_logic.v(17691)
  // ../RTL/cortexm0ds_logic.v(19991)
  // ../RTL/cortexm0ds_logic.v(18291)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~(D*B)*~(~C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0011001011111010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6_reg  (
    .a({_al_u4081_o,open_n77892}),
    .b({_al_u4191_o,open_n77893}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xs1iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/K84iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I74iu6 }),
    .f({_al_u5767_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tkdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Acebx6 }));  // ../RTL/cortexm0ds_logic.v(19991)
  // ../RTL/cortexm0ds_logic.v(18211)
  // ../RTL/cortexm0ds_logic.v(18199)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 ,open_n77908}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ws4iu6_lutinv ,open_n77909}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dg2qw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx8ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eg7iu6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T24iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/O34iu6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .f({_al_u5663_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xf7iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tyaax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2bax6 }));  // ../RTL/cortexm0ds_logic.v(18211)
  // ../RTL/cortexm0ds_logic.v(18738)
  // ../RTL/cortexm0ds_logic.v(20003)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("~(C*B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1111111100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tzebx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eclax6_reg  (
    .b({_al_u6958_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sjqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uvliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hfkiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6844_o,_al_u1910_o}),
    .mi({open_n77939,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zuliu6 ,_al_u1911_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r10_o[2] }));  // ../RTL/cortexm0ds_logic.v(18738)
  // ../RTL/cortexm0ds_logic.v(18833)
  // ../RTL/cortexm0ds_logic.v(18841)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U0rax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vkqax6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[29] }));  // ../RTL/cortexm0ds_logic.v(18833)
  // ../RTL/cortexm0ds_logic.v(18832)
  // ../RTL/cortexm0ds_logic.v(18842)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U2rax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Viqax6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rimiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1liu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[27] }));  // ../RTL/cortexm0ds_logic.v(18832)
  // ../RTL/cortexm0ds_logic.v(19936)
  // ../RTL/cortexm0ds_logic.v(18326)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(~(~D*~B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0101111101001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6_reg  (
    .a({_al_u4061_o,_al_u1968_o}),
    .b({_al_u4225_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G64iu6 }),
    .f({_al_u5795_o,_al_u2173_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U4fax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hpbbx6 }));  // ../RTL/cortexm0ds_logic.v(19936)
  // ../RTL/cortexm0ds_logic.v(19641)
  // ../RTL/cortexm0ds_logic.v(19635)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gz6ax6 ,open_n78012}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1wpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpgiu6 ),
    .clk(XTAL1_wire),
    .d({_al_u6333_o,_al_u546_o}),
    .mi(\u_cmsdk_mcu/HWDATA [31:30]),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/prst_reg ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rerow6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mpgiu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uj4bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tl4bx6 }));  // ../RTL/cortexm0ds_logic.v(19641)
  // ../RTL/cortexm0ds_logic.v(18372)
  // ../RTL/cortexm0ds_logic.v(18366)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    //.LUTG0("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D)"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101001011100),
    .INIT_LUTF1(16'b0000111110101100),
    .INIT_LUTG0(16'b0000101001011100),
    .INIT_LUTG1(16'b0000111110101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6_reg  (
    .a({_al_u4490_o,_al_u4490_o}),
    .b({_al_u4537_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 }),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uofax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sqfax6 }));  // ../RTL/cortexm0ds_logic.v(18372)
  // ../RTL/cortexm0ds_logic.v(19995)
  // ../RTL/cortexm0ds_logic.v(20095)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~((C*~A)*~(D)*~(B)+(C*~A)*D*~(B)+~((C*~A))*D*B+(C*~A)*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001111101111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0010001111101111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6_reg  (
    .a({open_n78048,_al_u1253_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,_al_u1676_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1720_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kadbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bcdbx6 }),
    .f({_al_u1721_o,_al_u1718_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Urgbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ojebx6 }));  // ../RTL/cortexm0ds_logic.v(19995)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Usqax6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ickiu6 ),
    .clk(XTAL1_wire),
    .mi({open_n78078,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 }),
    .q({open_n78096,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r2_o[20] }));  // ../RTL/cortexm0ds_logic.v(18837)
  // ../RTL/cortexm0ds_logic.v(18908)
  // ../RTL/cortexm0ds_logic.v(18914)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V1vax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wpuax6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C7miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4liu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[29] }));  // ../RTL/cortexm0ds_logic.v(18908)
  // ../RTL/cortexm0ds_logic.v(18910)
  // ../RTL/cortexm0ds_logic.v(18916)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V5vax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vtuax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Voqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r1_o[25] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Admiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hsliu6 }),
    .f({_al_u1247_o,_al_u1196_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[16] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[25] }));  // ../RTL/cortexm0ds_logic.v(18910)
  // ../RTL/cortexm0ds_logic.v(18911)
  // ../RTL/cortexm0ds_logic.v(18918)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V9vax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vvuax6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jlmiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fyliu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[21] }));  // ../RTL/cortexm0ds_logic.v(18911)
  // ../RTL/cortexm0ds_logic.v(18903)
  // ../RTL/cortexm0ds_logic.v(18919)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vbvax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yfuax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[6] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bomiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Sokiu6 }),
    .f({_al_u1095_o,_al_u1113_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[12] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[6] }));  // ../RTL/cortexm0ds_logic.v(18903)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vltpw6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .mi({open_n78184,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qcaiu6 }),
    .q({open_n78202,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[2] }));  // ../RTL/cortexm0ds_logic.v(17687)
  // ../RTL/cortexm0ds_logic.v(18913)
  // ../RTL/cortexm0ds_logic.v(18912)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vxuax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vzuax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[19] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E1miu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D4miu6 }),
    .f({_al_u1163_o,_al_u1154_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[20] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[19] }));  // ../RTL/cortexm0ds_logic.v(18913)
  // ../RTL/cortexm0ds_logic.v(18298)
  // ../RTL/cortexm0ds_logic.v(19966)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6_reg  (
    .a({_al_u4035_o,open_n78221}),
    .b({_al_u4101_o,open_n78222}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ns8ax6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Td7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y84iu6 ,open_n78226}),
    .f({_al_u5764_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X44iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W0dbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yxdax6 }));  // ../RTL/cortexm0ds_logic.v(18298)
  // ../RTL/cortexm0ds_logic.v(18315)
  // ../RTL/cortexm0ds_logic.v(19950)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*~A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000101110111011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6_reg  (
    .a({_al_u4071_o,_al_u1925_o}),
    .b({_al_u4096_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lcqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ae7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R84iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U64iu6 }),
    .f({_al_u5789_o,_al_u2210_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wfcbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gkeax6 }));  // ../RTL/cortexm0ds_logic.v(18315)
  // ../RTL/cortexm0ds_logic.v(18915)
  // ../RTL/cortexm0ds_logic.v(18909)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wruax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V3vax6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Eqqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kmqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r7_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r6_o[17] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wckiu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uoliu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 }),
    .f({_al_u1145_o,_al_u1137_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[1] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r4_o[17] }));  // ../RTL/cortexm0ds_logic.v(18915)
  // ../RTL/cortexm0ds_logic.v(19977)
  // ../RTL/cortexm0ds_logic.v(18164)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*~A))"),
    //.LUTF1("(~(C*~B)*~(D*~A))"),
    //.LUTG0("(~(D*C)*~(B*~A))"),
    //.LUTG1("(~(C*~B)*~(D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101110111011),
    .INIT_LUTF1(16'b1000101011001111),
    .INIT_LUTG0(16'b0000101110111011),
    .INIT_LUTG1(16'b1000101011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I3lhu6 ,_al_u2225_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y5lhu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Gdqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zg7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wvgax6 }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N64iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B74iu6 }),
    .f({_al_u5481_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qoyow6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xc9ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fldbx6 }));  // ../RTL/cortexm0ds_logic.v(19977)
  // ../RTL/cortexm0ds_logic.v(18251)
  // ../RTL/cortexm0ds_logic.v(18258)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("((D@B)*(C@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001001001001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6_reg  (
    .a({_al_u4056_o,open_n78292}),
    .b({_al_u4219_o,open_n78293}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/He7iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Iqzhu6_lutinv }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oh4iu6 ,open_n78304}),
    .f({_al_u5754_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z54iu6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xdcax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0cax6 }));  // ../RTL/cortexm0ds_logic.v(18251)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xkqpw6_reg  (
    .c({open_n78313,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Utqpw6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n267 ),
    .clk(SWCLKTCK_pad),
    .d({open_n78314,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qwfax6 }),
    .mi({open_n78325,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cjqpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kxhpw6 ),
    .f({open_n78326,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n267 }),
    .q({open_n78330,\u_cmsdk_mcu/u_cmsdk_mcu_system/cpu0cdbgpwrupreq }));  // ../RTL/cortexm0ds_logic.v(17572)
  // ../RTL/cortexm0ds_logic.v(18016)
  // ../RTL/cortexm0ds_logic.v(18007)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C*~D))"),
    //.LUT1("~(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001111110011),
    .INIT_LUT1(16'b1100000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6_reg  (
    .b({_al_u5053_o,_al_u5830_o}),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Df4iu6 }),
    .clk(XTAL1_wire),
    .d({_al_u5349_o,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/n382 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xu2qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 }));  // ../RTL/cortexm0ds_logic.v(18016)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6_reg  (
    .clk(XTAL1_wire),
    .mi({open_n78371,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xvqpw6 }),
    .sr(\u_cmsdk_mcu/u_cmsdk_mcu_clkctrl/dbgrst_reg ),
    .q({open_n78377,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xxqpw6 }));  // ../RTL/cortexm0ds_logic.v(17593)
  // ../RTL/cortexm0ds_logic.v(19784)
  // ../RTL/cortexm0ds_logic.v(17703)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7upw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zr7bx6_reg  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Cpqow6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Fnqow6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[15] }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Lf8iu6 ),
    .clk(XTAL1_wire),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r5_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] }),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bamiu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .f({_al_u1138_o,_al_u1132_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r0_o[15] }));  // ../RTL/cortexm0ds_logic.v(19784)
  // ../RTL/cortexm0ds_logic.v(19975)
  // ../RTL/cortexm0ds_logic.v(17817)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6_reg  (
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xl1iu6_lutinv }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 }),
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C53iu6 ),
    .clk(SWCLKTCK_pad),
    .d({_al_u1703_o,_al_u1712_o}),
    .mi({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Hlwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Jfdbx6 }),
    .f({_al_u1704_o,_al_u1713_o}),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ymwpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ahdbx6 }));  // ../RTL/cortexm0ds_logic.v(19975)
  // ../RTL/cortexm0ds_logic.v(17964)
  // ../RTL/cortexm0ds_logic.v(17479)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~A*~(D*B))"),
    //.LUTF1("~(C*~A*~(D*B))"),
    //.LUTG0("~(C*~A*~(D*B))"),
    //.LUTG1("~(C*~A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110111110101111),
    .INIT_LUTF1(16'b1110111110101111),
    .INIT_LUTG0(16'b1110111110101111),
    .INIT_LUTG1(16'b1110111110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6_reg|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6_reg  (
    .a({_al_u1743_o,_al_u1743_o}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vk1iu6 }),
    .c({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ay1iu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S02iu6 }),
    .clk(SWCLKTCK_pad),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uunpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X42qw6 }),
    .q({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zwnpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C72qw6 }));  // ../RTL/cortexm0ds_logic.v(17964)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zx7bx6_reg  (
    .ce(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pckiu6 ),
    .clk(XTAL1_wire),
    .mi({open_n78457,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zfmiu6 }),
    .q({open_n78464,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_r3_o[15] }));  // ../RTL/cortexm0ds_logic.v(19787)
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qehbx6 ,1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E4yhu6 ,open_n78465}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [1],open_n78485}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u1  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xn7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vj3qw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dugax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ksgax6 }),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [3:2]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u4|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u3  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pg3qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P23qw6 }),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c3 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [5:4]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u6|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u5  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vn9bx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Bf3qw6 }),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c5 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [7:6]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u8|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u7  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ke1qw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nd3qw6 }),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c7 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [9:8]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/u9_al_u7279  (
    .a({open_n78578,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Yf1qw6 }),
    .b({open_n78579,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add0/c9 ),
    .f({open_n78598,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrkbx6 [10]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u11_al_u7251  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c11 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [11]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c15 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u15_al_u7252  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c15 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [17],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [15]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c19 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u19_al_u7253  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c19 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [21],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [19]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c23 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [22],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u23_al_u7254  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c23 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [25],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [23]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c27 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [26],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u27_al_u7255  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c27 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [29],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [27]}),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [30],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u3_al_u7249  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c3 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [3]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c7 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/u7_al_u7250  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c7 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [7]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c11 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/ucin_al_u7248  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[1] ,1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[0] }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [1],open_n78748}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add1/c3 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Zsfpw6 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u11_al_u7259  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[14] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[12] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[15] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[13] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c11 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [12]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c15 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [13]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u15_al_u7260  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[18] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[16] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[19] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[17] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c15 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [16]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c19 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [19],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [17]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u19_al_u7261  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[22] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[20] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[23] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[21] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c19 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [22],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [20]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c23 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [23],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [21]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u23_al_u7262  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[26] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[24] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[27] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[25] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c23 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [26],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [24]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c27 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [27],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [25]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u27_al_u7263  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[30] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[28] }),
    .b({open_n78823,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[29] }),
    .c(2'b00),
    .d(2'b00),
    .e({open_n78826,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c27 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [30],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [28]}),
    .fx({open_n78842,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [29]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u3_al_u7257  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[6] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[4] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[7] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[5] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c3 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [4]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c7 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [5]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/u7_al_u7258  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[10] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[8] }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[11] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[9] }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c7 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [8]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c11 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [9]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/ucin_al_u7256  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[2] ,1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/vis_pc_o[3] ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/R0ghu6 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [2],open_n78898}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add2/c3 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N5fpw6 [3],open_n78899}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u11_al_u7242  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q1epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/C1epw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X1epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/J1epw6 }),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [11]}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [12]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c11 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [12]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c15 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [15],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [13]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u15_al_u7243  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/G3epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L2epw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N3epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z2epw6 }),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [17],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [15]}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [16]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c15 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [16]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c19 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [19],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [17]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u19_al_u7244  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/I4epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/U3epw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P4epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/B4epw6 }),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [21],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [19]}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [22],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [20]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c19 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [22],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [20]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c23 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [23],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [21]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u23_al_u7245  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [25],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [23]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [26],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [24]}),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [25],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [23]}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [26],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [24]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c23 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [26],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [24]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c27 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [27],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [25]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u27_al_u7246  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [29],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [27]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [30],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [28]}),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [29],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [27]}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [30],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [28]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c27 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [30],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [28]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c31 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [31],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [29]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u31_al_u7247  (
    .a({open_n78992,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/D5epw6 }),
    .c(2'b00),
    .d({open_n78997,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [31]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c31 ),
    .f({open_n79014,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [32]}),
    .fx({open_n79016,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [33]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u3_al_u7240  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [3]}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/E2epw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [4]}),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [3]}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [4]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c3 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [4]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c7 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [7],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [5]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/u7_al_u7241  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Q5phu6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/S2epw6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/W4epw6 }),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [7]}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [8]}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c7 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [8]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c11 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [11],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [9]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/ucin_al_u7239  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [1],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Dqfhu6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Qbfpw6 [0]}),
    .c(2'b00),
    .d({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [1],1'b1}),
    .e({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Idfpw6 [0]}),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [2],open_n79072}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add3_u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/add4/c3 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [3],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nxkbx6 [1]}));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [17:0]),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [17:0]),
    .p({open_n79158,open_n79159,open_n79160,open_n79161,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_31 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_30 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_29 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_28 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_27 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_26 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_25 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_24 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_23 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_22 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_21 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_20 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_19 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_18 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_17 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_16 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_15 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_14 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_0_0 }));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [17:0]),
    .b({4'b0000,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [31:18]}),
    .p({open_n79245,open_n79246,open_n79247,open_n79248,open_n79249,open_n79250,open_n79251,open_n79252,open_n79253,open_n79254,open_n79255,open_n79256,open_n79257,open_n79258,open_n79259,open_n79260,open_n79261,open_n79262,open_n79263,open_n79264,open_n79265,open_n79266,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_0_1_0 }));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_  (
    .a({4'b0000,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Mifpw6 [31:18]}),
    .b(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tgfpw6 [17:0]),
    .p({open_n79350,open_n79351,open_n79352,open_n79353,open_n79354,open_n79355,open_n79356,open_n79357,open_n79358,open_n79359,open_n79360,open_n79361,open_n79362,open_n79363,open_n79364,open_n79365,open_n79366,open_n79367,open_n79368,open_n79369,open_n79370,open_n79371,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_13 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_12 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_11 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_10 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_9 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_8 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_7 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_5 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_4 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_3 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_2 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_1 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/mult0_1_0_0 }));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u11_al_u7267  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/T9kpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Pt7ax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rfxax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/V0jpw6 }),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c11 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [13],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [11]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c15 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [14],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u15_al_u7268  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Amupw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nbxax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N0xpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Wlspw6 }),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c15 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [17],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [15]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c19 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [18],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u19_al_u7269  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Tjkpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Nr7ax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/F9gbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Z8jpw6 }),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c19 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [21],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [19]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c23 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [22],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u23_al_u7270  (
    .a({open_n79426,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Coupw6 }),
    .c(2'b11),
    .d({open_n79431,1'b0}),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c23 ),
    .f({open_n79448,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [23]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u3_al_u7265  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Y7opw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/P0ibx6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Rv7ax6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Johbx6 }),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c3 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [5],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [3]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c7 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [6],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/u7_al_u7266  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Uojbx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ujxax6 }),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vrtpw6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Ss0qw6 }),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c7 ),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [9],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [7]}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c11 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [10],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/ucin_al_u7264  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Oarpw6 ,1'b0}),
    .b({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Kzabx6 ,\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/N8rpw6 }),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [1],open_n79507}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub0/c3 ),
    .fx({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [2],\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/L6gpw6 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/ucin  (
    .a({\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/X5phu6 ,1'b0}),
    .b({1'b1,open_n79510}),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u2|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u1  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [1:0]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c1 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [2:1]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u4|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u3  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [3:2]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c3 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [4:3]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u6|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u5  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [5:4]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c5 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [6:5]),
    .fco(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u0|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u8|u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/u7  (
    .a(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Vnfpw6 [7:6]),
    .b(2'b00),
    .fci(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/sub1/c7 ),
    .f(\u_cmsdk_mcu/u_cmsdk_mcu_system/u_cortex_m0_integration/u_logic/Xlfpw6 [8:7]));

endmodule 

